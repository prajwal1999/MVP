-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity dotP_even is -- 
  generic (tag_length : integer); 
  port ( -- 
    R : in  std_logic_vector(7 downto 0);
    result : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity dotP_even;
architecture dotP_even_arch of dotP_even is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal R_buffer :  std_logic_vector(7 downto 0);
  signal R_update_enable: Boolean;
  -- output port buffer signals
  signal result_buffer :  std_logic_vector(31 downto 0);
  signal result_update_enable: Boolean;
  signal dotP_even_CP_0_start: Boolean;
  signal dotP_even_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_20_branch_ack_0 : boolean;
  signal do_while_stmt_20_branch_req_0 : boolean;
  signal phi_stmt_22_req_1 : boolean;
  signal phi_stmt_22_req_0 : boolean;
  signal phi_stmt_22_ack_0 : boolean;
  signal nC_153_26_buf_req_0 : boolean;
  signal nC_153_26_buf_ack_0 : boolean;
  signal nC_153_26_buf_req_1 : boolean;
  signal nC_153_26_buf_ack_1 : boolean;
  signal phi_stmt_27_req_1 : boolean;
  signal phi_stmt_27_req_0 : boolean;
  signal phi_stmt_27_ack_0 : boolean;
  signal nval_0_98_31_buf_req_0 : boolean;
  signal nval_0_98_31_buf_ack_0 : boolean;
  signal nval_0_98_31_buf_req_1 : boolean;
  signal nval_0_98_31_buf_ack_1 : boolean;
  signal phi_stmt_32_req_1 : boolean;
  signal phi_stmt_32_req_0 : boolean;
  signal phi_stmt_32_ack_0 : boolean;
  signal nval_1_113_36_buf_req_0 : boolean;
  signal nval_1_113_36_buf_ack_0 : boolean;
  signal nval_1_113_36_buf_req_1 : boolean;
  signal nval_1_113_36_buf_ack_1 : boolean;
  signal phi_stmt_37_req_1 : boolean;
  signal phi_stmt_37_req_0 : boolean;
  signal phi_stmt_37_ack_0 : boolean;
  signal nval_2_128_41_buf_req_0 : boolean;
  signal nval_2_128_41_buf_ack_0 : boolean;
  signal nval_2_128_41_buf_req_1 : boolean;
  signal nval_2_128_41_buf_ack_1 : boolean;
  signal phi_stmt_42_req_1 : boolean;
  signal phi_stmt_42_req_0 : boolean;
  signal phi_stmt_42_ack_0 : boolean;
  signal array_obj_ref_71_load_0_req_0 : boolean;
  signal array_obj_ref_71_load_0_ack_0 : boolean;
  signal nval_3_143_46_buf_req_0 : boolean;
  signal nval_3_143_46_buf_ack_0 : boolean;
  signal nval_3_143_46_buf_req_1 : boolean;
  signal nval_3_143_46_buf_ack_1 : boolean;
  signal array_obj_ref_56_index_0_scale_req_0 : boolean;
  signal array_obj_ref_56_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_56_index_0_scale_req_1 : boolean;
  signal array_obj_ref_56_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_56_index_sum_1_req_0 : boolean;
  signal array_obj_ref_56_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_56_index_sum_1_req_1 : boolean;
  signal array_obj_ref_56_index_sum_1_ack_1 : boolean;
  signal ADD_u32_u32_167_inst_ack_1 : boolean;
  signal array_obj_ref_56_load_0_req_0 : boolean;
  signal array_obj_ref_56_load_0_ack_0 : boolean;
  signal ADD_u8_u8_152_inst_ack_1 : boolean;
  signal array_obj_ref_56_load_0_req_1 : boolean;
  signal array_obj_ref_56_load_0_ack_1 : boolean;
  signal ADD_u32_u32_167_inst_req_1 : boolean;
  signal ADD_u8_u8_152_inst_req_1 : boolean;
  signal array_obj_ref_61_index_0_scale_req_0 : boolean;
  signal array_obj_ref_61_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_61_index_0_scale_req_1 : boolean;
  signal array_obj_ref_61_index_0_scale_ack_1 : boolean;
  signal ADD_u8_u8_152_inst_ack_0 : boolean;
  signal array_obj_ref_61_index_sum_1_req_0 : boolean;
  signal array_obj_ref_61_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_61_index_sum_1_req_1 : boolean;
  signal array_obj_ref_61_index_sum_1_ack_1 : boolean;
  signal ADD_u32_u32_167_inst_ack_0 : boolean;
  signal ADD_u32_u32_167_inst_req_0 : boolean;
  signal ADD_u8_u8_152_inst_req_0 : boolean;
  signal array_obj_ref_61_load_0_req_0 : boolean;
  signal array_obj_ref_61_load_0_ack_0 : boolean;
  signal array_obj_ref_61_load_0_req_1 : boolean;
  signal array_obj_ref_61_load_0_ack_1 : boolean;
  signal array_obj_ref_66_index_0_scale_req_0 : boolean;
  signal array_obj_ref_66_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_66_index_0_scale_req_1 : boolean;
  signal array_obj_ref_66_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_66_index_sum_1_req_0 : boolean;
  signal array_obj_ref_66_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_66_index_sum_1_req_1 : boolean;
  signal array_obj_ref_66_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_66_load_0_req_0 : boolean;
  signal array_obj_ref_66_load_0_ack_0 : boolean;
  signal W_val_3_126_delayed_5_0_134_inst_ack_1 : boolean;
  signal array_obj_ref_66_load_0_req_1 : boolean;
  signal array_obj_ref_66_load_0_ack_1 : boolean;
  signal do_while_stmt_20_branch_ack_1 : boolean;
  signal W_val_3_126_delayed_5_0_134_inst_req_1 : boolean;
  signal array_obj_ref_71_index_0_scale_req_0 : boolean;
  signal array_obj_ref_71_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_71_index_0_scale_req_1 : boolean;
  signal array_obj_ref_71_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_71_index_sum_1_req_0 : boolean;
  signal array_obj_ref_71_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_71_index_sum_1_req_1 : boolean;
  signal array_obj_ref_71_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_71_load_0_req_1 : boolean;
  signal array_obj_ref_71_load_0_ack_1 : boolean;
  signal array_obj_ref_75_load_0_req_0 : boolean;
  signal array_obj_ref_75_load_0_ack_0 : boolean;
  signal array_obj_ref_75_load_0_req_1 : boolean;
  signal array_obj_ref_75_load_0_ack_1 : boolean;
  signal array_obj_ref_79_load_0_req_0 : boolean;
  signal array_obj_ref_79_load_0_ack_0 : boolean;
  signal array_obj_ref_79_load_0_req_1 : boolean;
  signal array_obj_ref_79_load_0_ack_1 : boolean;
  signal array_obj_ref_83_load_0_req_0 : boolean;
  signal array_obj_ref_83_load_0_ack_0 : boolean;
  signal array_obj_ref_83_load_0_req_1 : boolean;
  signal array_obj_ref_83_load_0_ack_1 : boolean;
  signal array_obj_ref_87_load_0_req_0 : boolean;
  signal array_obj_ref_87_load_0_ack_0 : boolean;
  signal array_obj_ref_87_load_0_req_1 : boolean;
  signal array_obj_ref_87_load_0_ack_1 : boolean;
  signal W_val_0_90_delayed_5_0_89_inst_req_0 : boolean;
  signal W_val_0_90_delayed_5_0_89_inst_ack_0 : boolean;
  signal W_val_0_90_delayed_5_0_89_inst_req_1 : boolean;
  signal W_val_0_90_delayed_5_0_89_inst_ack_1 : boolean;
  signal W_val_1_102_delayed_5_0_104_inst_req_0 : boolean;
  signal W_val_1_102_delayed_5_0_104_inst_ack_0 : boolean;
  signal W_val_1_102_delayed_5_0_104_inst_req_1 : boolean;
  signal W_val_1_102_delayed_5_0_104_inst_ack_1 : boolean;
  signal W_val_2_114_delayed_5_0_119_inst_req_0 : boolean;
  signal W_val_2_114_delayed_5_0_119_inst_ack_0 : boolean;
  signal W_val_2_114_delayed_5_0_119_inst_req_1 : boolean;
  signal W_val_2_114_delayed_5_0_119_inst_ack_1 : boolean;
  signal W_val_3_126_delayed_5_0_134_inst_req_0 : boolean;
  signal W_val_3_126_delayed_5_0_134_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "dotP_even_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 8) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= R;
  R_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(tag_length + 7 downto 8) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 7 downto 8);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  dotP_even_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "dotP_even_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= result_buffer;
  result <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= dotP_even_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= dotP_even_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= dotP_even_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  dotP_even_CP_0: Block -- control-path 
    signal dotP_even_CP_0_elements: BooleanArray(202 downto 0);
    -- 
  begin -- 
    dotP_even_CP_0_elements(0) <= dotP_even_CP_0_start;
    dotP_even_CP_0_symbol <= dotP_even_CP_0_elements(202);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_19/$entry
      -- CP-element group 0: 	 branch_block_stmt_19/branch_block_stmt_19__entry__
      -- CP-element group 0: 	 branch_block_stmt_19/do_while_stmt_20__entry__
      -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	200 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	202 
    -- CP-element group 1: 	201 
    -- CP-element group 1:  members (10) 
      -- CP-element group 1: 	 branch_block_stmt_19/$exit
      -- CP-element group 1: 	 branch_block_stmt_19/branch_block_stmt_19__exit__
      -- CP-element group 1: 	 branch_block_stmt_19/do_while_stmt_20__exit__
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_Update/cr
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_Update/$entry
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_Sample/rr
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_update_start_
      -- CP-element group 1: 	 assign_stmt_168/ADD_u32_u32_167_sample_start_
      -- CP-element group 1: 	 assign_stmt_168/$entry
      -- 
    cr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(1), ack => ADD_u32_u32_167_inst_req_1); -- 
    rr_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(1), ack => ADD_u32_u32_167_inst_req_0); -- 
    dotP_even_CP_0_elements(1) <= dotP_even_CP_0_elements(200);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_19/do_while_stmt_20/$entry
      -- CP-element group 2: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20__entry__
      -- 
    dotP_even_CP_0_elements(2) <= dotP_even_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	200 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20__exit__
      -- 
    -- Element group dotP_even_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_19/do_while_stmt_20/loop_back
      -- 
    -- Element group dotP_even_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	198 
    -- CP-element group 5: 	199 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/condition_done
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/$entry
      -- 
    dotP_even_CP_0_elements(5) <= dotP_even_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	197 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_19/do_while_stmt_20/loop_body_done
      -- 
    dotP_even_CP_0_elements(6) <= dotP_even_CP_0_elements(197);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	95 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/back_edge_to_loop_body
      -- 
    dotP_even_CP_0_elements(7) <= dotP_even_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	97 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/first_time_through_loop_body
      -- 
    dotP_even_CP_0_elements(8) <= dotP_even_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	112 
    -- CP-element group 9: 	116 
    -- CP-element group 9: 	124 
    -- CP-element group 9: 	125 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	196 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	151 
    -- CP-element group 9: 	142 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	90 
    -- CP-element group 9: 	111 
    -- CP-element group 9:  members (26) 
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_0/index_resize_ack
      -- 
    -- Element group dotP_even_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	195 
    -- CP-element group 10: 	196 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/condition_evaluated
      -- 
    condition_evaluated_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(10), ack => do_while_stmt_20_branch_req_0); -- 
    dotP_even_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(14) & dotP_even_CP_0_elements(195) & dotP_even_CP_0_elements(196);
      gj_dotP_even_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	89 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	91 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_start__ps
      -- 
    dotP_even_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(15) & dotP_even_CP_0_elements(32) & dotP_even_CP_0_elements(51) & dotP_even_CP_0_elements(70) & dotP_even_CP_0_elements(89) & dotP_even_CP_0_elements(14);
      gj_dotP_even_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	92 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	122 
    -- CP-element group 12: 	181 
    -- CP-element group 12: 	185 
    -- CP-element group 12: 	189 
    -- CP-element group 12: 	177 
    -- CP-element group 12: 	173 
    -- CP-element group 12: 	169 
    -- CP-element group 12: 	193 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	161 
    -- CP-element group 12: 	148 
    -- CP-element group 12: 	165 
    -- CP-element group 12: 	109 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	89 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_sample_completed_
      -- 
    dotP_even_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(17) & dotP_even_CP_0_elements(35) & dotP_even_CP_0_elements(54) & dotP_even_CP_0_elements(73) & dotP_even_CP_0_elements(92);
      gj_dotP_even_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	90 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	93 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_start__ps
      -- 
    dotP_even_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(16) & dotP_even_CP_0_elements(33) & dotP_even_CP_0_elements(52) & dotP_even_CP_0_elements(71) & dotP_even_CP_0_elements(90);
      gj_dotP_even_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	94 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/aggregated_phi_update_ack
      -- 
    dotP_even_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(37) & dotP_even_CP_0_elements(56) & dotP_even_CP_0_elements(75) & dotP_even_CP_0_elements(94);
      gj_dotP_even_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	195 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_start_
      -- 
    dotP_even_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(195);
      gj_dotP_even_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	130 
    -- CP-element group 16: 	174 
    -- CP-element group 16: 	170 
    -- CP-element group 16: 	194 
    -- CP-element group 16: 	166 
    -- CP-element group 16: 	156 
    -- CP-element group 16: 	162 
    -- CP-element group 16: 	143 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_start_
      -- 
    dotP_even_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 1,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1,8 => 0,9 => 1);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(117) & dotP_even_CP_0_elements(130) & dotP_even_CP_0_elements(174) & dotP_even_CP_0_elements(170) & dotP_even_CP_0_elements(194) & dotP_even_CP_0_elements(166) & dotP_even_CP_0_elements(156) & dotP_even_CP_0_elements(162) & dotP_even_CP_0_elements(143);
      gj_dotP_even_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_sample_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	115 
    -- CP-element group 18: 	128 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	172 
    -- CP-element group 18: 	168 
    -- CP-element group 18: 	192 
    -- CP-element group 18: 	160 
    -- CP-element group 18: 	154 
    -- CP-element group 18: 	164 
    -- CP-element group 18: 	141 
    -- CP-element group 18:  members (150) 
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_word_addrgen/root_register_ack
      -- 
    -- Element group dotP_even_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_trigger
      -- 
    dotP_even_CP_0_elements(19) <= dotP_even_CP_0_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_loopback_sample_req_ps
      -- 
    phi_stmt_22_loopback_sample_req_39_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_22_loopback_sample_req_39_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(20), ack => phi_stmt_22_req_1); -- 
    -- Element group dotP_even_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_trigger
      -- 
    dotP_even_CP_0_elements(21) <= dotP_even_CP_0_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_entry_sample_req_ps
      -- 
    phi_stmt_22_entry_sample_req_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_22_entry_sample_req_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(22), ack => phi_stmt_22_req_0); -- 
    -- Element group dotP_even_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_22_phi_mux_ack_ps
      -- 
    phi_stmt_22_phi_mux_ack_45_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_22_ack_0, ack => dotP_even_CP_0_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_sample_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_start_
      -- 
    -- Element group dotP_even_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_completed__ps
      -- 
    dotP_even_CP_0_elements(26) <= dotP_even_CP_0_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_25_update_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(25), ack => dotP_even_CP_0_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Sample/req
      -- 
    req_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(28), ack => nC_153_26_buf_req_0); -- 
    -- Element group dotP_even_CP_0_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_update_start_
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Update/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(29), ack => nC_153_26_buf_req_1); -- 
    -- Element group dotP_even_CP_0_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Sample/ack
      -- 
    ack_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nC_153_26_buf_ack_0, ack => dotP_even_CP_0_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nC_26_Update/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nC_153_26_buf_ack_1, ack => dotP_even_CP_0_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	120 
    -- CP-element group 32: 	12 
    -- CP-element group 32: 	179 
    -- CP-element group 32: 	163 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_sample_start_
      -- 
    dotP_even_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(120) & dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(179) & dotP_even_CP_0_elements(163);
      gj_dotP_even_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	178 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_update_start_
      -- 
    dotP_even_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(178);
      gj_dotP_even_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_sample_start__ps
      -- 
    dotP_even_CP_0_elements(34) <= dotP_even_CP_0_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_sample_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_update_start__ps
      -- 
    dotP_even_CP_0_elements(36) <= dotP_even_CP_0_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	176 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_update_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_loopback_trigger
      -- 
    dotP_even_CP_0_elements(38) <= dotP_even_CP_0_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_loopback_sample_req_ps
      -- 
    phi_stmt_27_loopback_sample_req_83_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_27_loopback_sample_req_83_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(39), ack => phi_stmt_27_req_1); -- 
    -- Element group dotP_even_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_entry_trigger
      -- 
    dotP_even_CP_0_elements(40) <= dotP_even_CP_0_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_entry_sample_req_ps
      -- 
    phi_stmt_27_entry_sample_req_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_27_entry_sample_req_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(41), ack => phi_stmt_27_req_0); -- 
    -- Element group dotP_even_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_27_phi_mux_ack_ps
      -- 
    phi_stmt_27_phi_mux_ack_89_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_27_ack_0, ack => dotP_even_CP_0_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_sample_start__ps
      -- 
    -- Element group dotP_even_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_update_start_
      -- 
    -- Element group dotP_even_CP_0_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_update_completed__ps
      -- 
    dotP_even_CP_0_elements(45) <= dotP_even_CP_0_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_30_update_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(44), ack => dotP_even_CP_0_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Sample/req
      -- 
    req_110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(47), ack => nval_0_98_31_buf_req_0); -- 
    -- Element group dotP_even_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_update_start_
      -- CP-element group 48: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Update/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(48), ack => nval_0_98_31_buf_req_1); -- 
    -- Element group dotP_even_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Sample/ack
      -- 
    ack_111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_0_98_31_buf_ack_0, ack => dotP_even_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_0_31_Update/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_0_98_31_buf_ack_1, ack => dotP_even_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: 	183 
    -- CP-element group 51: 	167 
    -- CP-element group 51: 	133 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_sample_start_
      -- 
    dotP_even_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(183) & dotP_even_CP_0_elements(167) & dotP_even_CP_0_elements(133);
      gj_dotP_even_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	182 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_update_start_
      -- 
    dotP_even_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(182);
      gj_dotP_even_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_sample_start__ps
      -- 
    dotP_even_CP_0_elements(53) <= dotP_even_CP_0_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_sample_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_update_start__ps
      -- 
    dotP_even_CP_0_elements(55) <= dotP_even_CP_0_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	180 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_update_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_loopback_trigger
      -- 
    dotP_even_CP_0_elements(57) <= dotP_even_CP_0_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_loopback_sample_req_ps
      -- 
    phi_stmt_32_loopback_sample_req_127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_32_loopback_sample_req_127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(58), ack => phi_stmt_32_req_1); -- 
    -- Element group dotP_even_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_entry_trigger
      -- 
    dotP_even_CP_0_elements(59) <= dotP_even_CP_0_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_entry_sample_req_ps
      -- 
    phi_stmt_32_entry_sample_req_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_32_entry_sample_req_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(60), ack => phi_stmt_32_req_0); -- 
    -- Element group dotP_even_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_32_phi_mux_ack_ps
      -- 
    phi_stmt_32_phi_mux_ack_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_32_ack_0, ack => dotP_even_CP_0_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_sample_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_update_start_
      -- 
    -- Element group dotP_even_CP_0_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_update_completed__ps
      -- 
    dotP_even_CP_0_elements(64) <= dotP_even_CP_0_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_35_update_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(63), ack => dotP_even_CP_0_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Sample/req
      -- 
    req_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(66), ack => nval_1_113_36_buf_req_0); -- 
    -- Element group dotP_even_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_update_start_
      -- CP-element group 67: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Update/req
      -- 
    req_159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(67), ack => nval_1_113_36_buf_req_1); -- 
    -- Element group dotP_even_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Sample/ack
      -- 
    ack_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_1_113_36_buf_ack_0, ack => dotP_even_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_1_36_Update/ack
      -- 
    ack_160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_1_113_36_buf_ack_1, ack => dotP_even_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	187 
    -- CP-element group 70: 	171 
    -- CP-element group 70: 	146 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_sample_start_
      -- 
    dotP_even_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(187) & dotP_even_CP_0_elements(171) & dotP_even_CP_0_elements(146);
      gj_dotP_even_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	186 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_update_start_
      -- 
    dotP_even_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(186);
      gj_dotP_even_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_sample_start__ps
      -- 
    dotP_even_CP_0_elements(72) <= dotP_even_CP_0_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_sample_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_update_start__ps
      -- 
    dotP_even_CP_0_elements(74) <= dotP_even_CP_0_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	184 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_update_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_loopback_trigger
      -- 
    dotP_even_CP_0_elements(76) <= dotP_even_CP_0_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_loopback_sample_req_ps
      -- 
    phi_stmt_37_loopback_sample_req_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_37_loopback_sample_req_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(77), ack => phi_stmt_37_req_1); -- 
    -- Element group dotP_even_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_entry_trigger
      -- 
    dotP_even_CP_0_elements(78) <= dotP_even_CP_0_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_entry_sample_req_ps
      -- 
    phi_stmt_37_entry_sample_req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_37_entry_sample_req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(79), ack => phi_stmt_37_req_0); -- 
    -- Element group dotP_even_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_37_phi_mux_ack
      -- 
    phi_stmt_37_phi_mux_ack_177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_37_ack_0, ack => dotP_even_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_sample_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_update_start_
      -- 
    -- Element group dotP_even_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_update_completed__ps
      -- 
    dotP_even_CP_0_elements(83) <= dotP_even_CP_0_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_40_update_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(82), ack => dotP_even_CP_0_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Sample/req
      -- 
    req_198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(85), ack => nval_2_128_41_buf_req_0); -- 
    -- Element group dotP_even_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_update_start_
      -- CP-element group 86: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Update/req
      -- 
    req_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(86), ack => nval_2_128_41_buf_req_1); -- 
    -- Element group dotP_even_CP_0_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Sample/ack
      -- 
    ack_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_2_128_41_buf_ack_0, ack => dotP_even_CP_0_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_2_41_Update/ack
      -- 
    ack_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_2_128_41_buf_ack_1, ack => dotP_even_CP_0_elements(88)); -- 
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	12 
    -- CP-element group 89: 	175 
    -- CP-element group 89: 	191 
    -- CP-element group 89: 	159 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	11 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_sample_start_
      -- 
    dotP_even_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(175) & dotP_even_CP_0_elements(191) & dotP_even_CP_0_elements(159);
      gj_dotP_even_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	9 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	190 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	13 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_update_start_
      -- 
    dotP_even_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_even_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(190);
      gj_dotP_even_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	11 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_sample_start__ps
      -- 
    dotP_even_CP_0_elements(91) <= dotP_even_CP_0_elements(11);
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	12 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_sample_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(92) is bound as output of CP function.
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	13 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_update_start__ps
      -- 
    dotP_even_CP_0_elements(93) <= dotP_even_CP_0_elements(13);
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: 	188 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_update_completed__ps
      -- 
    -- Element group dotP_even_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	7 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_loopback_trigger
      -- 
    dotP_even_CP_0_elements(95) <= dotP_even_CP_0_elements(7);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_loopback_sample_req
      -- CP-element group 96: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_loopback_sample_req_ps
      -- 
    phi_stmt_42_loopback_sample_req_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_42_loopback_sample_req_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(96), ack => phi_stmt_42_req_1); -- 
    -- Element group dotP_even_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	8 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_entry_trigger
      -- 
    dotP_even_CP_0_elements(97) <= dotP_even_CP_0_elements(8);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_entry_sample_req
      -- CP-element group 98: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_entry_sample_req_ps
      -- 
    phi_stmt_42_entry_sample_req_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_42_entry_sample_req_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(98), ack => phi_stmt_42_req_0); -- 
    -- Element group dotP_even_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_phi_mux_ack
      -- CP-element group 99: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/phi_stmt_42_phi_mux_ack_ps
      -- 
    phi_stmt_42_phi_mux_ack_221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_42_ack_0, ack => dotP_even_CP_0_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_sample_completed__ps
      -- CP-element group 100: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_sample_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_update_start_
      -- 
    -- Element group dotP_even_CP_0_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_update_completed__ps
      -- 
    dotP_even_CP_0_elements(102) <= dotP_even_CP_0_elements(103);
    -- CP-element group 103:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	102 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/type_cast_45_update_completed_
      -- 
    -- Element group dotP_even_CP_0_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(101), ack => dotP_even_CP_0_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Sample/req
      -- 
    req_242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(104), ack => nval_3_143_46_buf_req_0); -- 
    -- Element group dotP_even_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_update_start_
      -- CP-element group 105: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Update/req
      -- 
    req_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(105), ack => nval_3_143_46_buf_req_1); -- 
    -- Element group dotP_even_CP_0_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Sample/ack
      -- 
    ack_243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_3_143_46_buf_ack_0, ack => dotP_even_CP_0_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/R_nval_3_46_Update/ack
      -- 
    ack_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_3_143_46_buf_ack_1, ack => dotP_even_CP_0_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	118 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	119 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/word_0/rr
      -- 
    rr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(108), ack => array_obj_ref_56_load_0_req_0); -- 
    dotP_even_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(118) & dotP_even_CP_0_elements(119);
      gj_dotP_even_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	12 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	120 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	120 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_update_start_
      -- CP-element group 109: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/$entry
      -- CP-element group 109: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/word_0/cr
      -- 
    cr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(109), ack => array_obj_ref_56_load_0_req_1); -- 
    dotP_even_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(120);
      gj_dotP_even_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	114 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	117 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	115 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scaled_0
      -- 
    dotP_even_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(114) & dotP_even_CP_0_elements(117);
      gj_dotP_even_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_sample_start
      -- CP-element group 111: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Sample/rr
      -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(111), ack => array_obj_ref_56_index_0_scale_req_0); -- 
    dotP_even_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(113);
      gj_dotP_even_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	9 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_update_start
      -- CP-element group 112: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Update/cr
      -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(112), ack => array_obj_ref_56_index_0_scale_req_1); -- 
    dotP_even_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(114);
      gj_dotP_even_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	197 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_sample_complete
      -- CP-element group 113: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Sample/ra
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_index_0_scale_ack_0, ack => dotP_even_CP_0_elements(113)); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	110 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_update_complete
      -- CP-element group 114: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_index_scale_0_Update/ca
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_index_0_scale_ack_1, ack => dotP_even_CP_0_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	18 
    -- CP-element group 115: 	110 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_sample_start
      -- CP-element group 115: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Sample/rr
      -- 
    rr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(115), ack => array_obj_ref_56_index_sum_1_req_0); -- 
    dotP_even_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(110) & dotP_even_CP_0_elements(117);
      gj_dotP_even_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	119 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_update_start
      -- CP-element group 116: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Update/cr
      -- 
    cr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(116), ack => array_obj_ref_56_index_sum_1_req_1); -- 
    dotP_even_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(119);
      gj_dotP_even_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	197 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	16 
    -- CP-element group 117: 	110 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_sample_complete
      -- CP-element group 117: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Sample/ra
      -- 
    ra_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_index_sum_1_ack_0, ack => dotP_even_CP_0_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	108 
    -- CP-element group 118:  members (18) 
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_word_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_root_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_offset_calculated
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_update_complete
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_partial_sum_1_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_final_index_sum_regn/$entry
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_final_index_sum_regn/$exit
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_final_index_sum_regn/req
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_final_index_sum_regn/ack
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_base_plus_offset/$entry
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_base_plus_offset/$exit
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_base_plus_offset/sum_rename_req
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_base_plus_offset/sum_rename_ack
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_word_addrgen/$entry
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_word_addrgen/$exit
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_word_addrgen/root_register_req
      -- CP-element group 118: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_word_addrgen/root_register_ack
      -- 
    ca_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_index_sum_1_ack_1, ack => dotP_even_CP_0_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: 	108 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Sample/word_access_start/word_0/ra
      -- 
    ra_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_load_0_ack_0, ack => dotP_even_CP_0_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	109 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	197 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	32 
    -- CP-element group 120: 	109 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/array_obj_ref_56_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/array_obj_ref_56_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/array_obj_ref_56_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_56_Update/array_obj_ref_56_Merge/merge_ack
      -- 
    ca_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_56_load_0_ack_1, ack => dotP_even_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	131 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	132 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	132 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/$entry
      -- CP-element group 121: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/word_0/$entry
      -- CP-element group 121: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/word_0/rr
      -- 
    rr_430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(121), ack => array_obj_ref_61_load_0_req_0); -- 
    dotP_even_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(131) & dotP_even_CP_0_elements(132);
      gj_dotP_even_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	12 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	133 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	133 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_update_start_
      -- CP-element group 122: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/$entry
      -- CP-element group 122: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/word_0/$entry
      -- CP-element group 122: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/word_0/cr
      -- 
    cr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(122), ack => array_obj_ref_61_load_0_req_1); -- 
    dotP_even_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(133);
      gj_dotP_even_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	130 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scaled_0
      -- 
    dotP_even_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(127) & dotP_even_CP_0_elements(130);
      gj_dotP_even_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	9 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_sample_start
      -- CP-element group 124: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Sample/rr
      -- 
    rr_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(124), ack => array_obj_ref_61_index_0_scale_req_0); -- 
    dotP_even_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(126);
      gj_dotP_even_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	9 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_update_start
      -- CP-element group 125: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Update/cr
      -- 
    cr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(125), ack => array_obj_ref_61_index_0_scale_req_1); -- 
    dotP_even_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(127);
      gj_dotP_even_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	197 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Sample/ra
      -- 
    ra_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_0_scale_ack_0, ack => dotP_even_CP_0_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_update_complete
      -- CP-element group 127: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_index_scale_0_Update/ca
      -- 
    ca_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_0_scale_ack_1, ack => dotP_even_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	18 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_sample_start
      -- CP-element group 128: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Sample/rr
      -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(128), ack => array_obj_ref_61_index_sum_1_req_0); -- 
    dotP_even_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(123) & dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(130);
      gj_dotP_even_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	132 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_update_start
      -- CP-element group 129: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Update/cr
      -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(129), ack => array_obj_ref_61_index_sum_1_req_1); -- 
    dotP_even_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(132);
      gj_dotP_even_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	197 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	123 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	16 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_sample_complete
      -- CP-element group 130: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_sum_1_ack_0, ack => dotP_even_CP_0_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	121 
    -- CP-element group 131:  members (18) 
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_word_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_root_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_offset_calculated
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_update_complete
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_partial_sum_1_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_final_index_sum_regn/$entry
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_final_index_sum_regn/$exit
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_final_index_sum_regn/req
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_final_index_sum_regn/ack
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_base_plus_offset/$entry
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_base_plus_offset/$exit
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_base_plus_offset/sum_rename_req
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_base_plus_offset/sum_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_word_addrgen/$entry
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_word_addrgen/$exit
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_word_addrgen/root_register_req
      -- CP-element group 131: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_word_addrgen/root_register_ack
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_sum_1_ack_1, ack => dotP_even_CP_0_elements(131)); -- 
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	121 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	121 
    -- CP-element group 132: 	129 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/$exit
      -- CP-element group 132: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/word_0/$exit
      -- CP-element group 132: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Sample/word_access_start/word_0/ra
      -- 
    ra_431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_load_0_ack_0, ack => dotP_even_CP_0_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	122 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	197 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	122 
    -- CP-element group 133: 	51 
    -- CP-element group 133:  members (9) 
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/$exit
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/word_0/$exit
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/word_access_complete/word_0/ca
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/array_obj_ref_61_Merge/$entry
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/array_obj_ref_61_Merge/$exit
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/array_obj_ref_61_Merge/merge_req
      -- CP-element group 133: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_61_Update/array_obj_ref_61_Merge/merge_ack
      -- 
    ca_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_load_0_ack_1, ack => dotP_even_CP_0_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	144 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	145 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	145 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/$entry
      -- CP-element group 134: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/word_0/rr
      -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(134), ack => array_obj_ref_66_load_0_req_0); -- 
    dotP_even_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(144) & dotP_even_CP_0_elements(145);
      gj_dotP_even_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	146 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	146 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_update_start_
      -- CP-element group 135: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/$entry
      -- CP-element group 135: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 135: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/word_0/cr
      -- 
    cr_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(135), ack => array_obj_ref_66_load_0_req_1); -- 
    dotP_even_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(146);
      gj_dotP_even_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	140 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	143 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scaled_0
      -- 
    dotP_even_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(140) & dotP_even_CP_0_elements(143);
      gj_dotP_even_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_sample_start
      -- CP-element group 137: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Sample/rr
      -- 
    rr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(137), ack => array_obj_ref_66_index_0_scale_req_0); -- 
    dotP_even_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(139);
      gj_dotP_even_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_update_start
      -- CP-element group 138: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Update/cr
      -- 
    cr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(138), ack => array_obj_ref_66_index_0_scale_req_1); -- 
    dotP_even_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(140);
      gj_dotP_even_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	197 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_sample_complete
      -- CP-element group 139: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Sample/ra
      -- 
    ra_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_index_0_scale_ack_0, ack => dotP_even_CP_0_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	136 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_update_complete
      -- CP-element group 140: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_index_scale_0_Update/ca
      -- 
    ca_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_index_0_scale_ack_1, ack => dotP_even_CP_0_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	18 
    -- CP-element group 141: 	136 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_sample_start
      -- CP-element group 141: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Sample/rr
      -- 
    rr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(141), ack => array_obj_ref_66_index_sum_1_req_0); -- 
    dotP_even_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(136) & dotP_even_CP_0_elements(143);
      gj_dotP_even_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	9 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	145 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_update_start
      -- CP-element group 142: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Update/cr
      -- 
    cr_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(142), ack => array_obj_ref_66_index_sum_1_req_1); -- 
    dotP_even_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(145);
      gj_dotP_even_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	197 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	16 
    -- CP-element group 143: 	136 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_sample_complete
      -- CP-element group 143: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Sample/ra
      -- 
    ra_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_index_sum_1_ack_0, ack => dotP_even_CP_0_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	134 
    -- CP-element group 144:  members (18) 
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_root_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_offset_calculated
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_word_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_update_complete
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_partial_sum_1_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_final_index_sum_regn/$entry
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_final_index_sum_regn/$exit
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_final_index_sum_regn/req
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_final_index_sum_regn/ack
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_base_plus_offset/$entry
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_base_plus_offset/$exit
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_base_plus_offset/sum_rename_req
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_word_addrgen/$entry
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_word_addrgen/$exit
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_word_addrgen/root_register_req
      -- CP-element group 144: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_word_addrgen/root_register_ack
      -- 
    ca_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_index_sum_1_ack_1, ack => dotP_even_CP_0_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	134 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	134 
    -- CP-element group 145: 	142 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Sample/word_access_start/word_0/ra
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_load_0_ack_0, ack => dotP_even_CP_0_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	135 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	197 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	135 
    -- CP-element group 146: 	70 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/array_obj_ref_66_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/array_obj_ref_66_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/array_obj_ref_66_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_66_Update/array_obj_ref_66_Merge/merge_ack
      -- 
    ca_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_66_load_0_ack_1, ack => dotP_even_CP_0_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	157 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	158 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	158 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/$entry
      -- CP-element group 147: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/word_0/$entry
      -- CP-element group 147: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/word_0/rr
      -- CP-element group 147: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_sample_start_
      -- 
    rr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(147), ack => array_obj_ref_71_load_0_req_0); -- 
    dotP_even_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(157) & dotP_even_CP_0_elements(158);
      gj_dotP_even_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	12 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	159 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	159 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/$entry
      -- CP-element group 148: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/word_0/$entry
      -- CP-element group 148: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_update_start_
      -- CP-element group 148: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/word_0/cr
      -- 
    cr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(148), ack => array_obj_ref_71_load_0_req_1); -- 
    dotP_even_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(159);
      gj_dotP_even_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	153 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	156 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scaled_0
      -- 
    dotP_even_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(153) & dotP_even_CP_0_elements(156);
      gj_dotP_even_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_sample_start
      -- CP-element group 150: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Sample/rr
      -- 
    rr_570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(150), ack => array_obj_ref_71_index_0_scale_req_0); -- 
    dotP_even_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(152);
      gj_dotP_even_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	9 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_update_start
      -- CP-element group 151: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Update/cr
      -- 
    cr_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(151), ack => array_obj_ref_71_index_0_scale_req_1); -- 
    dotP_even_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(153);
      gj_dotP_even_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	197 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_sample_complete
      -- CP-element group 152: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Sample/ra
      -- 
    ra_571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_0_scale_ack_0, ack => dotP_even_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	149 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_update_complete
      -- CP-element group 153: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_index_scale_0_Update/ca
      -- 
    ca_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_0_scale_ack_1, ack => dotP_even_CP_0_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	18 
    -- CP-element group 154: 	149 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_sample_start
      -- CP-element group 154: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Sample/rr
      -- 
    rr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(154), ack => array_obj_ref_71_index_sum_1_req_0); -- 
    dotP_even_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(149) & dotP_even_CP_0_elements(156);
      gj_dotP_even_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	158 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_update_start
      -- CP-element group 155: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Update/cr
      -- 
    cr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(155), ack => array_obj_ref_71_index_sum_1_req_1); -- 
    dotP_even_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(9) & dotP_even_CP_0_elements(158);
      gj_dotP_even_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	197 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	16 
    -- CP-element group 156: 	154 
    -- CP-element group 156: 	149 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_sample_complete
      -- CP-element group 156: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Sample/ra
      -- 
    ra_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_sum_1_ack_0, ack => dotP_even_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	147 
    -- CP-element group 157:  members (18) 
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_final_index_sum_regn/$entry
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_final_index_sum_regn/$exit
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_final_index_sum_regn/req
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_final_index_sum_regn/ack
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_base_plus_offset/$entry
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_base_plus_offset/$exit
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_base_plus_offset/sum_rename_req
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_base_plus_offset/sum_rename_ack
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_word_addrgen/$entry
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_word_addrgen/$exit
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_word_addrgen/root_register_req
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_word_addrgen/root_register_ack
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_word_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_root_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_offset_calculated
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_update_complete
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_partial_sum_1_Update/ca
      -- 
    ca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_sum_1_ack_1, ack => dotP_even_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	147 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: 	147 
    -- CP-element group 158:  members (5) 
      -- CP-element group 158: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/$exit
      -- CP-element group 158: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Sample/word_access_start/word_0/ra
      -- CP-element group 158: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_sample_completed_
      -- 
    ra_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_load_0_ack_0, ack => dotP_even_CP_0_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	148 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	197 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	148 
    -- CP-element group 159: 	89 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/$exit
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/word_0/$exit
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/word_access_complete/word_0/ca
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/array_obj_ref_71_Merge/$entry
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/array_obj_ref_71_Merge/$exit
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/array_obj_ref_71_Merge/merge_req
      -- CP-element group 159: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_71_Update/array_obj_ref_71_Merge/merge_ack
      -- 
    ca_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_load_0_ack_1, ack => dotP_even_CP_0_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	18 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/$entry
      -- CP-element group 160: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/word_0/rr
      -- 
    rr_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(160), ack => array_obj_ref_75_load_0_req_0); -- 
    dotP_even_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(162);
      gj_dotP_even_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	12 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_update_start_
      -- CP-element group 161: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/$entry
      -- CP-element group 161: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/word_0/cr
      -- 
    cr_702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(161), ack => array_obj_ref_75_load_0_req_1); -- 
    dotP_even_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(163);
      gj_dotP_even_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	16 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Sample/word_access_start/word_0/ra
      -- 
    ra_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_load_0_ack_0, ack => dotP_even_CP_0_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	197 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	32 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/array_obj_ref_75_Merge/$entry
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/array_obj_ref_75_Merge/$exit
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/array_obj_ref_75_Merge/merge_req
      -- CP-element group 163: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_75_Update/array_obj_ref_75_Merge/merge_ack
      -- 
    ca_703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_load_0_ack_1, ack => dotP_even_CP_0_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	18 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/$entry
      -- CP-element group 164: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/word_0/$entry
      -- CP-element group 164: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/word_0/rr
      -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(164), ack => array_obj_ref_79_load_0_req_0); -- 
    dotP_even_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(166);
      gj_dotP_even_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	12 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_update_start_
      -- CP-element group 165: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/$entry
      -- CP-element group 165: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/word_0/$entry
      -- CP-element group 165: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/word_0/cr
      -- 
    cr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(165), ack => array_obj_ref_79_load_0_req_1); -- 
    dotP_even_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(167);
      gj_dotP_even_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	16 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/$exit
      -- CP-element group 166: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/word_0/$exit
      -- CP-element group 166: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Sample/word_access_start/word_0/ra
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_79_load_0_ack_0, ack => dotP_even_CP_0_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	197 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: 	51 
    -- CP-element group 167:  members (9) 
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/$exit
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/word_0/$exit
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/word_access_complete/word_0/ca
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/array_obj_ref_79_Merge/$entry
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/array_obj_ref_79_Merge/$exit
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/array_obj_ref_79_Merge/merge_req
      -- CP-element group 167: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_79_Update/array_obj_ref_79_Merge/merge_ack
      -- 
    ca_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_79_load_0_ack_1, ack => dotP_even_CP_0_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	18 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/$entry
      -- CP-element group 168: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/word_0/rr
      -- 
    rr_817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(168), ack => array_obj_ref_83_load_0_req_0); -- 
    dotP_even_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(170);
      gj_dotP_even_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	12 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_update_start_
      -- CP-element group 169: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/$entry
      -- CP-element group 169: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/word_0/$entry
      -- CP-element group 169: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/word_0/cr
      -- 
    cr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(169), ack => array_obj_ref_83_load_0_req_1); -- 
    dotP_even_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(171);
      gj_dotP_even_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	16 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (5) 
      -- CP-element group 170: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/$exit
      -- CP-element group 170: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/word_0/$exit
      -- CP-element group 170: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Sample/word_access_start/word_0/ra
      -- 
    ra_818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_83_load_0_ack_0, ack => dotP_even_CP_0_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	197 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	70 
    -- CP-element group 171:  members (9) 
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/$exit
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/word_0/$exit
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/word_access_complete/word_0/ca
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/array_obj_ref_83_Merge/$entry
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/array_obj_ref_83_Merge/$exit
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/array_obj_ref_83_Merge/merge_req
      -- CP-element group 171: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_83_Update/array_obj_ref_83_Merge/merge_ack
      -- 
    ca_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_83_load_0_ack_1, ack => dotP_even_CP_0_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	18 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (5) 
      -- CP-element group 172: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/$entry
      -- CP-element group 172: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/word_0/rr
      -- 
    rr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(172), ack => array_obj_ref_87_load_0_req_0); -- 
    dotP_even_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(174);
      gj_dotP_even_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	12 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_update_start_
      -- CP-element group 173: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/$entry
      -- CP-element group 173: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/word_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/word_0/cr
      -- 
    cr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(173), ack => array_obj_ref_87_load_0_req_1); -- 
    dotP_even_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(175);
      gj_dotP_even_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	16 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/$exit
      -- CP-element group 174: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/word_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Sample/word_access_start/word_0/ra
      -- 
    ra_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_87_load_0_ack_0, ack => dotP_even_CP_0_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	197 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	89 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/$exit
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/word_0/$exit
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/word_access_complete/word_0/ca
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/array_obj_ref_87_Merge/$entry
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/array_obj_ref_87_Merge/$exit
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/array_obj_ref_87_Merge/merge_req
      -- CP-element group 175: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/array_obj_ref_87_Update/array_obj_ref_87_Merge/merge_ack
      -- 
    ca_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_87_load_0_ack_1, ack => dotP_even_CP_0_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	37 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Sample/req
      -- 
    req_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(176), ack => W_val_0_90_delayed_5_0_89_inst_req_0); -- 
    dotP_even_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(37) & dotP_even_CP_0_elements(178);
      gj_dotP_even_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	12 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_update_start_
      -- CP-element group 177: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Update/req
      -- 
    req_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(177), ack => W_val_0_90_delayed_5_0_89_inst_req_1); -- 
    dotP_even_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(179);
      gj_dotP_even_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	33 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Sample/ack
      -- 
    ack_906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_0_90_delayed_5_0_89_inst_ack_0, ack => dotP_even_CP_0_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	197 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	32 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_91_Update/ack
      -- 
    ack_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_0_90_delayed_5_0_89_inst_ack_1, ack => dotP_even_CP_0_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	56 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Sample/req
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(180), ack => W_val_1_102_delayed_5_0_104_inst_req_0); -- 
    dotP_even_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(56) & dotP_even_CP_0_elements(182);
      gj_dotP_even_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	12 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_update_start_
      -- CP-element group 181: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Update/req
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(181), ack => W_val_1_102_delayed_5_0_104_inst_req_1); -- 
    dotP_even_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(183);
      gj_dotP_even_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	52 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Sample/ack
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_1_102_delayed_5_0_104_inst_ack_0, ack => dotP_even_CP_0_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	197 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: 	51 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_106_Update/ack
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_1_102_delayed_5_0_104_inst_ack_1, ack => dotP_even_CP_0_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	75 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Sample/req
      -- 
    req_933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(184), ack => W_val_2_114_delayed_5_0_119_inst_req_0); -- 
    dotP_even_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(75) & dotP_even_CP_0_elements(186);
      gj_dotP_even_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	12 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_update_start_
      -- CP-element group 185: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Update/req
      -- 
    req_938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(185), ack => W_val_2_114_delayed_5_0_119_inst_req_1); -- 
    dotP_even_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(187);
      gj_dotP_even_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	71 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Sample/ack
      -- 
    ack_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_2_114_delayed_5_0_119_inst_ack_0, ack => dotP_even_CP_0_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	197 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	70 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_121_Update/ack
      -- 
    ack_939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_2_114_delayed_5_0_119_inst_ack_1, ack => dotP_even_CP_0_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	94 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Sample/req
      -- 
    req_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(188), ack => W_val_3_126_delayed_5_0_134_inst_req_0); -- 
    dotP_even_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(94) & dotP_even_CP_0_elements(190);
      gj_dotP_even_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	12 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Update/req
      -- CP-element group 189: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_update_start_
      -- 
    req_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(189), ack => W_val_3_126_delayed_5_0_134_inst_req_1); -- 
    dotP_even_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(191);
      gj_dotP_even_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: 	90 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Sample/ack
      -- 
    ack_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_3_126_delayed_5_0_134_inst_ack_0, ack => dotP_even_CP_0_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	197 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	89 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Update/ack
      -- CP-element group 191: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/assign_stmt_136_update_completed_
      -- 
    ack_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_3_126_delayed_5_0_134_inst_ack_1, ack => dotP_even_CP_0_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	18 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_sample_start_
      -- 
    rr_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(192), ack => ADD_u8_u8_152_inst_req_0); -- 
    dotP_even_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(18) & dotP_even_CP_0_elements(194);
      gj_dotP_even_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	12 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Update/cr
      -- CP-element group 193: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_update_start_
      -- 
    cr_966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_even_CP_0_elements(193), ack => ADD_u8_u8_152_inst_req_1); -- 
    dotP_even_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(12) & dotP_even_CP_0_elements(195);
      gj_dotP_even_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	16 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_sample_completed_
      -- 
    ra_962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_152_inst_ack_0, ack => dotP_even_CP_0_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	10 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	15 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/ADD_u8_u8_152_update_completed_
      -- 
    ca_967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_152_inst_ack_1, ack => dotP_even_CP_0_elements(195)); -- 
    -- CP-element group 196:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	9 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	10 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group dotP_even_CP_0_elements(196) is a control-delay.
    cp_element_196_delay: control_delay_element  generic map(name => " 196_delay", delay_value => 1)  port map(req => dotP_even_CP_0_elements(9), ack => dotP_even_CP_0_elements(196), clk => clk, reset =>reset);
    -- CP-element group 197:  join  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	117 
    -- CP-element group 197: 	113 
    -- CP-element group 197: 	120 
    -- CP-element group 197: 	126 
    -- CP-element group 197: 	130 
    -- CP-element group 197: 	183 
    -- CP-element group 197: 	187 
    -- CP-element group 197: 	175 
    -- CP-element group 197: 	179 
    -- CP-element group 197: 	171 
    -- CP-element group 197: 	191 
    -- CP-element group 197: 	167 
    -- CP-element group 197: 	133 
    -- CP-element group 197: 	139 
    -- CP-element group 197: 	159 
    -- CP-element group 197: 	152 
    -- CP-element group 197: 	156 
    -- CP-element group 197: 	146 
    -- CP-element group 197: 	163 
    -- CP-element group 197: 	143 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	6 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_19/do_while_stmt_20/do_while_stmt_20_loop_body/$exit
      -- 
    dotP_even_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 19) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15);
      constant place_markings: IntegerArray(0 to 19)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant place_delays: IntegerArray(0 to 19) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant joinName: string(1 to 30) := "dotP_even_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 20); -- 
    begin -- 
      preds <= dotP_even_CP_0_elements(117) & dotP_even_CP_0_elements(113) & dotP_even_CP_0_elements(120) & dotP_even_CP_0_elements(126) & dotP_even_CP_0_elements(130) & dotP_even_CP_0_elements(183) & dotP_even_CP_0_elements(187) & dotP_even_CP_0_elements(175) & dotP_even_CP_0_elements(179) & dotP_even_CP_0_elements(171) & dotP_even_CP_0_elements(191) & dotP_even_CP_0_elements(167) & dotP_even_CP_0_elements(133) & dotP_even_CP_0_elements(139) & dotP_even_CP_0_elements(159) & dotP_even_CP_0_elements(152) & dotP_even_CP_0_elements(156) & dotP_even_CP_0_elements(146) & dotP_even_CP_0_elements(163) & dotP_even_CP_0_elements(143);
      gj_dotP_even_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 20, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_even_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	5 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/ack
      -- CP-element group 198: 	 branch_block_stmt_19/do_while_stmt_20/loop_exit/$exit
      -- 
    ack_972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_20_branch_ack_0, ack => dotP_even_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	5 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/ack
      -- CP-element group 199: 	 branch_block_stmt_19/do_while_stmt_20/loop_taken/$exit
      -- 
    ack_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_20_branch_ack_1, ack => dotP_even_CP_0_elements(199)); -- 
    -- CP-element group 200:  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	3 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	1 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_19/do_while_stmt_20/$exit
      -- 
    dotP_even_CP_0_elements(200) <= dotP_even_CP_0_elements(3);
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	1 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_168/ADD_u32_u32_167_Sample/ra
      -- CP-element group 201: 	 assign_stmt_168/ADD_u32_u32_167_Sample/$exit
      -- CP-element group 201: 	 assign_stmt_168/ADD_u32_u32_167_sample_completed_
      -- 
    ra_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_167_inst_ack_0, ack => dotP_even_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	1 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (5) 
      -- CP-element group 202: 	 $exit
      -- CP-element group 202: 	 assign_stmt_168/ADD_u32_u32_167_Update/ca
      -- CP-element group 202: 	 assign_stmt_168/ADD_u32_u32_167_Update/$exit
      -- CP-element group 202: 	 assign_stmt_168/ADD_u32_u32_167_update_completed_
      -- CP-element group 202: 	 assign_stmt_168/$exit
      -- 
    ca_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_167_inst_ack_1, ack => dotP_even_CP_0_elements(202)); -- 
    dotP_even_do_while_stmt_20_terminator_977: loop_terminator -- 
      generic map (name => " dotP_even_do_while_stmt_20_terminator_977", max_iterations_in_flight =>15) 
      port map(loop_body_exit => dotP_even_CP_0_elements(6),loop_continue => dotP_even_CP_0_elements(199),loop_terminate => dotP_even_CP_0_elements(198),loop_back => dotP_even_CP_0_elements(4),loop_exit => dotP_even_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_22_phi_seq_73_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_even_CP_0_elements(21);
      dotP_even_CP_0_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_even_CP_0_elements(24);
      dotP_even_CP_0_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_even_CP_0_elements(26);
      dotP_even_CP_0_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_even_CP_0_elements(19);
      dotP_even_CP_0_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_even_CP_0_elements(30);
      dotP_even_CP_0_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_even_CP_0_elements(31);
      dotP_even_CP_0_elements(20) <= phi_mux_reqs(1);
      phi_stmt_22_phi_seq_73 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_22_phi_seq_73") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_even_CP_0_elements(11), 
          phi_sample_ack => dotP_even_CP_0_elements(17), 
          phi_update_req => dotP_even_CP_0_elements(13), 
          phi_update_ack => dotP_even_CP_0_elements(18), 
          phi_mux_ack => dotP_even_CP_0_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_27_phi_seq_117_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_even_CP_0_elements(40);
      dotP_even_CP_0_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_even_CP_0_elements(43);
      dotP_even_CP_0_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_even_CP_0_elements(45);
      dotP_even_CP_0_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_even_CP_0_elements(38);
      dotP_even_CP_0_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_even_CP_0_elements(49);
      dotP_even_CP_0_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_even_CP_0_elements(50);
      dotP_even_CP_0_elements(39) <= phi_mux_reqs(1);
      phi_stmt_27_phi_seq_117 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_27_phi_seq_117") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_even_CP_0_elements(34), 
          phi_sample_ack => dotP_even_CP_0_elements(35), 
          phi_update_req => dotP_even_CP_0_elements(36), 
          phi_update_ack => dotP_even_CP_0_elements(37), 
          phi_mux_ack => dotP_even_CP_0_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_32_phi_seq_161_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_even_CP_0_elements(59);
      dotP_even_CP_0_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_even_CP_0_elements(62);
      dotP_even_CP_0_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_even_CP_0_elements(64);
      dotP_even_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_even_CP_0_elements(57);
      dotP_even_CP_0_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_even_CP_0_elements(68);
      dotP_even_CP_0_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_even_CP_0_elements(69);
      dotP_even_CP_0_elements(58) <= phi_mux_reqs(1);
      phi_stmt_32_phi_seq_161 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_32_phi_seq_161") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_even_CP_0_elements(53), 
          phi_sample_ack => dotP_even_CP_0_elements(54), 
          phi_update_req => dotP_even_CP_0_elements(55), 
          phi_update_ack => dotP_even_CP_0_elements(56), 
          phi_mux_ack => dotP_even_CP_0_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_37_phi_seq_205_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_even_CP_0_elements(78);
      dotP_even_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_even_CP_0_elements(81);
      dotP_even_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_even_CP_0_elements(83);
      dotP_even_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_even_CP_0_elements(76);
      dotP_even_CP_0_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_even_CP_0_elements(87);
      dotP_even_CP_0_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_even_CP_0_elements(88);
      dotP_even_CP_0_elements(77) <= phi_mux_reqs(1);
      phi_stmt_37_phi_seq_205 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_37_phi_seq_205") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_even_CP_0_elements(72), 
          phi_sample_ack => dotP_even_CP_0_elements(73), 
          phi_update_req => dotP_even_CP_0_elements(74), 
          phi_update_ack => dotP_even_CP_0_elements(75), 
          phi_mux_ack => dotP_even_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_42_phi_seq_249_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_even_CP_0_elements(97);
      dotP_even_CP_0_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_even_CP_0_elements(100);
      dotP_even_CP_0_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_even_CP_0_elements(102);
      dotP_even_CP_0_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_even_CP_0_elements(95);
      dotP_even_CP_0_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_even_CP_0_elements(106);
      dotP_even_CP_0_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_even_CP_0_elements(107);
      dotP_even_CP_0_elements(96) <= phi_mux_reqs(1);
      phi_stmt_42_phi_seq_249 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_42_phi_seq_249") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_even_CP_0_elements(91), 
          phi_sample_ack => dotP_even_CP_0_elements(92), 
          phi_update_req => dotP_even_CP_0_elements(93), 
          phi_update_ack => dotP_even_CP_0_elements(94), 
          phi_mux_ack => dotP_even_CP_0_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_25_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= dotP_even_CP_0_elements(7);
        preds(1)  <= dotP_even_CP_0_elements(8);
        entry_tmerge_25 : transition_merge -- 
          generic map(name => " entry_tmerge_25")
          port map (preds => preds, symbol_out => dotP_even_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_165_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_166_wire : std_logic_vector(31 downto 0);
    signal C_22 : std_logic_vector(7 downto 0);
    signal Cr_52 : std_logic_vector(5 downto 0);
    signal MUL_u32_u32_111_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_126_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_141_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_96_wire : std_logic_vector(31 downto 0);
    signal R_Cr_55_resized : std_logic_vector(7 downto 0);
    signal R_Cr_55_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_60_resized : std_logic_vector(7 downto 0);
    signal R_Cr_60_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_65_resized : std_logic_vector(7 downto 0);
    signal R_Cr_65_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_70_resized : std_logic_vector(7 downto 0);
    signal R_Cr_70_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_74_resized : std_logic_vector(2 downto 0);
    signal R_Cr_74_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_78_resized : std_logic_vector(2 downto 0);
    signal R_Cr_78_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_82_resized : std_logic_vector(2 downto 0);
    signal R_Cr_82_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_86_resized : std_logic_vector(2 downto 0);
    signal R_Cr_86_scaled : std_logic_vector(2 downto 0);
    signal R_R_54_resized : std_logic_vector(7 downto 0);
    signal R_R_54_scaled : std_logic_vector(7 downto 0);
    signal R_R_59_resized : std_logic_vector(7 downto 0);
    signal R_R_59_scaled : std_logic_vector(7 downto 0);
    signal R_R_64_resized : std_logic_vector(7 downto 0);
    signal R_R_64_scaled : std_logic_vector(7 downto 0);
    signal R_R_69_resized : std_logic_vector(7 downto 0);
    signal R_R_69_scaled : std_logic_vector(7 downto 0);
    signal ULT_u8_u1_157_wire : std_logic_vector(0 downto 0);
    signal a_rc_0_57 : std_logic_vector(31 downto 0);
    signal a_rc_1_62 : std_logic_vector(31 downto 0);
    signal a_rc_2_67 : std_logic_vector(31 downto 0);
    signal a_rc_3_72 : std_logic_vector(31 downto 0);
    signal array_obj_ref_56_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_56_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_56_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_61_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_61_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_66_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_66_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_71_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_71_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_75_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_75_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_75_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_75_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_75_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_75_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_75_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_79_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_79_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_83_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_83_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_87_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_87_word_offset_0 : std_logic_vector(2 downto 0);
    signal konst_151_wire_constant : std_logic_vector(7 downto 0);
    signal konst_156_wire_constant : std_logic_vector(7 downto 0);
    signal nC_153 : std_logic_vector(7 downto 0);
    signal nC_153_26_buffered : std_logic_vector(7 downto 0);
    signal nval_0_98 : std_logic_vector(31 downto 0);
    signal nval_0_98_31_buffered : std_logic_vector(31 downto 0);
    signal nval_1_113 : std_logic_vector(31 downto 0);
    signal nval_1_113_36_buffered : std_logic_vector(31 downto 0);
    signal nval_2_128 : std_logic_vector(31 downto 0);
    signal nval_2_128_41_buffered : std_logic_vector(31 downto 0);
    signal nval_3_143 : std_logic_vector(31 downto 0);
    signal nval_3_143_46_buffered : std_logic_vector(31 downto 0);
    signal type_cast_25_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_30_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_35_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_40_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_45_wire_constant : std_logic_vector(31 downto 0);
    signal val_0_27 : std_logic_vector(31 downto 0);
    signal val_0_90_delayed_5_0_91 : std_logic_vector(31 downto 0);
    signal val_1_102_delayed_5_0_106 : std_logic_vector(31 downto 0);
    signal val_1_32 : std_logic_vector(31 downto 0);
    signal val_2_114_delayed_5_0_121 : std_logic_vector(31 downto 0);
    signal val_2_37 : std_logic_vector(31 downto 0);
    signal val_3_126_delayed_5_0_136 : std_logic_vector(31 downto 0);
    signal val_3_42 : std_logic_vector(31 downto 0);
    signal xval_0_76 : std_logic_vector(31 downto 0);
    signal xval_1_80 : std_logic_vector(31 downto 0);
    signal xval_2_84 : std_logic_vector(31 downto 0);
    signal xval_3_88 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_56_offset_scale_factor_0 <= "00001000";
    array_obj_ref_56_offset_scale_factor_1 <= "00000001";
    array_obj_ref_56_resized_base_address <= "00000000";
    array_obj_ref_56_word_offset_0 <= "00000000";
    array_obj_ref_61_offset_scale_factor_0 <= "00001000";
    array_obj_ref_61_offset_scale_factor_1 <= "00000001";
    array_obj_ref_61_resized_base_address <= "00000000";
    array_obj_ref_61_word_offset_0 <= "00000000";
    array_obj_ref_66_offset_scale_factor_0 <= "00001000";
    array_obj_ref_66_offset_scale_factor_1 <= "00000001";
    array_obj_ref_66_resized_base_address <= "00000000";
    array_obj_ref_66_word_offset_0 <= "00000000";
    array_obj_ref_71_offset_scale_factor_0 <= "00001000";
    array_obj_ref_71_offset_scale_factor_1 <= "00000001";
    array_obj_ref_71_resized_base_address <= "00000000";
    array_obj_ref_71_word_offset_0 <= "00000000";
    array_obj_ref_75_offset_scale_factor_0 <= "001";
    array_obj_ref_75_resized_base_address <= "000";
    array_obj_ref_75_word_offset_0 <= "000";
    array_obj_ref_79_offset_scale_factor_0 <= "001";
    array_obj_ref_79_resized_base_address <= "000";
    array_obj_ref_79_word_offset_0 <= "000";
    array_obj_ref_83_offset_scale_factor_0 <= "001";
    array_obj_ref_83_resized_base_address <= "000";
    array_obj_ref_83_word_offset_0 <= "000";
    array_obj_ref_87_offset_scale_factor_0 <= "001";
    array_obj_ref_87_resized_base_address <= "000";
    array_obj_ref_87_word_offset_0 <= "000";
    konst_151_wire_constant <= "00000100";
    konst_156_wire_constant <= "00100000";
    type_cast_25_wire_constant <= "00000000";
    type_cast_30_wire_constant <= "00000000000000000000000000000000";
    type_cast_35_wire_constant <= "00000000000000000000000000000000";
    type_cast_40_wire_constant <= "00000000000000000000000000000000";
    type_cast_45_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_22: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_25_wire_constant & nC_153_26_buffered;
      req <= phi_stmt_22_req_0 & phi_stmt_22_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_22",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_22_ack_0,
          idata => idata,
          odata => C_22,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_22
    phi_stmt_27: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_30_wire_constant & nval_0_98_31_buffered;
      req <= phi_stmt_27_req_0 & phi_stmt_27_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_27",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_27_ack_0,
          idata => idata,
          odata => val_0_27,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_27
    phi_stmt_32: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_35_wire_constant & nval_1_113_36_buffered;
      req <= phi_stmt_32_req_0 & phi_stmt_32_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_32",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_32_ack_0,
          idata => idata,
          odata => val_1_32,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_32
    phi_stmt_37: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_40_wire_constant & nval_2_128_41_buffered;
      req <= phi_stmt_37_req_0 & phi_stmt_37_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_37",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_37_ack_0,
          idata => idata,
          odata => val_2_37,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_37
    phi_stmt_42: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_45_wire_constant & nval_3_143_46_buffered;
      req <= phi_stmt_42_req_0 & phi_stmt_42_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_42",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_42_ack_0,
          idata => idata,
          odata => val_3_42,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_42
    -- flow-through slice operator slice_51_inst
    Cr_52 <= C_22(7 downto 2);
    W_val_0_90_delayed_5_0_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_0_90_delayed_5_0_89_inst_req_0;
      W_val_0_90_delayed_5_0_89_inst_ack_0<= wack(0);
      rreq(0) <= W_val_0_90_delayed_5_0_89_inst_req_1;
      W_val_0_90_delayed_5_0_89_inst_ack_1<= rack(0);
      W_val_0_90_delayed_5_0_89_inst : InterlockBuffer generic map ( -- 
        name => "W_val_0_90_delayed_5_0_89_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_0_27,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_0_90_delayed_5_0_91,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_1_102_delayed_5_0_104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_1_102_delayed_5_0_104_inst_req_0;
      W_val_1_102_delayed_5_0_104_inst_ack_0<= wack(0);
      rreq(0) <= W_val_1_102_delayed_5_0_104_inst_req_1;
      W_val_1_102_delayed_5_0_104_inst_ack_1<= rack(0);
      W_val_1_102_delayed_5_0_104_inst : InterlockBuffer generic map ( -- 
        name => "W_val_1_102_delayed_5_0_104_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_1_32,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_1_102_delayed_5_0_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_2_114_delayed_5_0_119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_2_114_delayed_5_0_119_inst_req_0;
      W_val_2_114_delayed_5_0_119_inst_ack_0<= wack(0);
      rreq(0) <= W_val_2_114_delayed_5_0_119_inst_req_1;
      W_val_2_114_delayed_5_0_119_inst_ack_1<= rack(0);
      W_val_2_114_delayed_5_0_119_inst : InterlockBuffer generic map ( -- 
        name => "W_val_2_114_delayed_5_0_119_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_2_37,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_2_114_delayed_5_0_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_3_126_delayed_5_0_134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_3_126_delayed_5_0_134_inst_req_0;
      W_val_3_126_delayed_5_0_134_inst_ack_0<= wack(0);
      rreq(0) <= W_val_3_126_delayed_5_0_134_inst_req_1;
      W_val_3_126_delayed_5_0_134_inst_ack_1<= rack(0);
      W_val_3_126_delayed_5_0_134_inst : InterlockBuffer generic map ( -- 
        name => "W_val_3_126_delayed_5_0_134_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_3_42,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_3_126_delayed_5_0_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nC_153_26_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nC_153_26_buf_req_0;
      nC_153_26_buf_ack_0<= wack(0);
      rreq(0) <= nC_153_26_buf_req_1;
      nC_153_26_buf_ack_1<= rack(0);
      nC_153_26_buf : InterlockBuffer generic map ( -- 
        name => "nC_153_26_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nC_153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nC_153_26_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_0_98_31_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_0_98_31_buf_req_0;
      nval_0_98_31_buf_ack_0<= wack(0);
      rreq(0) <= nval_0_98_31_buf_req_1;
      nval_0_98_31_buf_ack_1<= rack(0);
      nval_0_98_31_buf : InterlockBuffer generic map ( -- 
        name => "nval_0_98_31_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_0_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_0_98_31_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_1_113_36_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_1_113_36_buf_req_0;
      nval_1_113_36_buf_ack_0<= wack(0);
      rreq(0) <= nval_1_113_36_buf_req_1;
      nval_1_113_36_buf_ack_1<= rack(0);
      nval_1_113_36_buf : InterlockBuffer generic map ( -- 
        name => "nval_1_113_36_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_1_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_1_113_36_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_2_128_41_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_2_128_41_buf_req_0;
      nval_2_128_41_buf_ack_0<= wack(0);
      rreq(0) <= nval_2_128_41_buf_req_1;
      nval_2_128_41_buf_ack_1<= rack(0);
      nval_2_128_41_buf : InterlockBuffer generic map ( -- 
        name => "nval_2_128_41_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_2_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_2_128_41_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_3_143_46_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_3_143_46_buf_req_0;
      nval_3_143_46_buf_ack_0<= wack(0);
      rreq(0) <= nval_3_143_46_buf_req_1;
      nval_3_143_46_buf_ack_1<= rack(0);
      nval_3_143_46_buf : InterlockBuffer generic map ( -- 
        name => "nval_3_143_46_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_3_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_3_143_46_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_56_addr_0
    process(array_obj_ref_56_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_56_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_gather_scatter
    process(array_obj_ref_56_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_data_0;
      ov(31 downto 0) := iv;
      a_rc_0_57 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_54_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_index_1_rename
    process(R_Cr_55_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_55_resized;
      ov(7 downto 0) := iv;
      R_Cr_55_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_index_1_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov(5 downto 0) := iv;
      R_Cr_55_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_index_offset
    process(array_obj_ref_56_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_56_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_56_root_address_inst
    process(array_obj_ref_56_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_56_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_56_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_addr_0
    process(array_obj_ref_61_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_61_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_gather_scatter
    process(array_obj_ref_61_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_data_0;
      ov(31 downto 0) := iv;
      a_rc_1_62 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_59_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_rename
    process(R_Cr_60_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_60_resized;
      ov(7 downto 0) := iv;
      R_Cr_60_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov(5 downto 0) := iv;
      R_Cr_60_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_offset
    process(array_obj_ref_61_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_61_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_root_address_inst
    process(array_obj_ref_61_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_61_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_addr_0
    process(array_obj_ref_66_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_66_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_66_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_gather_scatter
    process(array_obj_ref_66_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_66_data_0;
      ov(31 downto 0) := iv;
      a_rc_2_67 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_64_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_index_1_rename
    process(R_Cr_65_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_65_resized;
      ov(7 downto 0) := iv;
      R_Cr_65_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_index_1_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov(5 downto 0) := iv;
      R_Cr_65_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_index_offset
    process(array_obj_ref_66_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_66_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_66_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_66_root_address_inst
    process(array_obj_ref_66_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_66_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_66_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_addr_0
    process(array_obj_ref_71_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_71_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_71_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_gather_scatter
    process(array_obj_ref_71_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_71_data_0;
      ov(31 downto 0) := iv;
      a_rc_3_72 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_69_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_index_1_rename
    process(R_Cr_70_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_70_resized;
      ov(7 downto 0) := iv;
      R_Cr_70_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_index_1_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov(5 downto 0) := iv;
      R_Cr_70_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_index_offset
    process(array_obj_ref_71_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_71_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_71_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_root_address_inst
    process(array_obj_ref_71_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_71_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_71_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_addr_0
    process(array_obj_ref_75_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_75_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_75_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_gather_scatter
    process(array_obj_ref_75_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_75_data_0;
      ov(31 downto 0) := iv;
      xval_0_76 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_0_rename
    process(R_Cr_74_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_74_resized;
      ov(2 downto 0) := iv;
      R_Cr_74_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_0_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov := iv(2 downto 0);
      R_Cr_74_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_offset
    process(R_Cr_74_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_74_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_75_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_root_address_inst
    process(array_obj_ref_75_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_75_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_75_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_addr_0
    process(array_obj_ref_79_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_79_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_79_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_gather_scatter
    process(array_obj_ref_79_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_79_data_0;
      ov(31 downto 0) := iv;
      xval_1_80 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_index_0_rename
    process(R_Cr_78_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_78_resized;
      ov(2 downto 0) := iv;
      R_Cr_78_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_index_0_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov := iv(2 downto 0);
      R_Cr_78_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_index_offset
    process(R_Cr_78_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_78_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_79_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_79_root_address_inst
    process(array_obj_ref_79_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_79_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_79_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_addr_0
    process(array_obj_ref_83_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_83_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_83_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_gather_scatter
    process(array_obj_ref_83_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_83_data_0;
      ov(31 downto 0) := iv;
      xval_2_84 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_index_0_rename
    process(R_Cr_82_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_82_resized;
      ov(2 downto 0) := iv;
      R_Cr_82_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_index_0_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov := iv(2 downto 0);
      R_Cr_82_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_index_offset
    process(R_Cr_82_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_82_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_83_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_83_root_address_inst
    process(array_obj_ref_83_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_83_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_83_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_addr_0
    process(array_obj_ref_87_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_87_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_87_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_gather_scatter
    process(array_obj_ref_87_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_87_data_0;
      ov(31 downto 0) := iv;
      xval_3_88 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_index_0_rename
    process(R_Cr_86_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_86_resized;
      ov(2 downto 0) := iv;
      R_Cr_86_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_index_0_resize
    process(Cr_52) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_52;
      ov := iv(2 downto 0);
      R_Cr_86_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_index_offset
    process(R_Cr_86_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_86_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_87_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_87_root_address_inst
    process(array_obj_ref_87_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_87_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_87_root_address <= ov(2 downto 0);
      --
    end process;
    do_while_stmt_20_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_157_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_20_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_20_branch_req_0,
          ack0 => do_while_stmt_20_branch_ack_0,
          ack1 => do_while_stmt_20_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_112_inst
    process(val_1_102_delayed_5_0_106, MUL_u32_u32_111_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_1_102_delayed_5_0_106, MUL_u32_u32_111_wire, tmp_var);
      nval_1_113 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_127_inst
    process(val_2_114_delayed_5_0_121, MUL_u32_u32_126_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_2_114_delayed_5_0_121, MUL_u32_u32_126_wire, tmp_var);
      nval_2_128 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_142_inst
    process(val_3_126_delayed_5_0_136, MUL_u32_u32_141_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_3_126_delayed_5_0_136, MUL_u32_u32_141_wire, tmp_var);
      nval_3_143 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_165_inst
    process(nval_2_128, nval_3_143) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nval_2_128, nval_3_143, tmp_var);
      ADD_u32_u32_165_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_166_inst
    process(nval_1_113, ADD_u32_u32_165_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nval_1_113, ADD_u32_u32_165_wire, tmp_var);
      ADD_u32_u32_166_wire <= tmp_var; --
    end process;
    -- shared split operator group (5) : ADD_u32_u32_167_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= nval_0_98 & ADD_u32_u32_166_wire;
      result_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_167_inst_req_0;
      ADD_u32_u32_167_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_167_inst_req_1;
      ADD_u32_u32_167_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_5_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- binary operator ADD_u32_u32_97_inst
    process(val_0_90_delayed_5_0_91, MUL_u32_u32_96_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_0_90_delayed_5_0_91, MUL_u32_u32_96_wire, tmp_var);
      nval_0_98 <= tmp_var; --
    end process;
    -- shared split operator group (7) : ADD_u8_u8_152_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= C_22;
      nC_153 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_152_inst_req_0;
      ADD_u8_u8_152_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_152_inst_req_1;
      ADD_u8_u8_152_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator MUL_u32_u32_111_inst
    process(a_rc_1_62, xval_1_80) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_1_62, xval_1_80, tmp_var);
      MUL_u32_u32_111_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_126_inst
    process(a_rc_2_67, xval_2_84) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_2_67, xval_2_84, tmp_var);
      MUL_u32_u32_126_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_141_inst
    process(a_rc_3_72, xval_3_88) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_3_72, xval_3_88, tmp_var);
      MUL_u32_u32_141_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_96_inst
    process(a_rc_0_57, xval_0_76) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_0_57, xval_0_76, tmp_var);
      MUL_u32_u32_96_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_157_inst
    process(nC_153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nC_153, konst_156_wire_constant, tmp_var);
      ULT_u8_u1_157_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_56_index_0_scale array_obj_ref_61_index_0_scale array_obj_ref_66_index_0_scale array_obj_ref_71_index_0_scale 
    ApIntMul_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      data_in <= R_R_54_resized & R_R_59_resized & R_R_64_resized & R_R_69_resized;
      R_R_54_scaled <= data_out(31 downto 24);
      R_R_59_scaled <= data_out(23 downto 16);
      R_R_64_scaled <= data_out(15 downto 8);
      R_R_69_scaled <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      reqL_unguarded(3) <= array_obj_ref_56_index_0_scale_req_0;
      reqL_unguarded(2) <= array_obj_ref_61_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_66_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_71_index_0_scale_req_0;
      array_obj_ref_56_index_0_scale_ack_0 <= ackL_unguarded(3);
      array_obj_ref_61_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_66_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_71_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_56_index_0_scale_req_1;
      reqR_unguarded(2) <= array_obj_ref_61_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_66_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_71_index_0_scale_req_1;
      array_obj_ref_56_index_0_scale_ack_1 <= ackR_unguarded(3);
      array_obj_ref_61_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_66_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_71_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_13_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_2: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_3: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_gI: SplitGuardInterface generic map(name => "ApIntMul_group_13_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_13",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00001000",
          constant_width => 8,
          use_constant  => true,
          full_rate  => true,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 4,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_56_index_sum_1 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_55_scaled & R_R_54_scaled;
      array_obj_ref_56_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_56_index_sum_1_req_0;
      array_obj_ref_56_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_56_index_sum_1_req_1;
      array_obj_ref_56_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_61_index_sum_1 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_60_scaled & R_R_59_scaled;
      array_obj_ref_61_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_61_index_sum_1_req_0;
      array_obj_ref_61_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_61_index_sum_1_req_1;
      array_obj_ref_61_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : array_obj_ref_66_index_sum_1 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_65_scaled & R_R_64_scaled;
      array_obj_ref_66_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_66_index_sum_1_req_0;
      array_obj_ref_66_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_66_index_sum_1_req_1;
      array_obj_ref_66_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : array_obj_ref_71_index_sum_1 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_70_scaled & R_R_69_scaled;
      array_obj_ref_71_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_71_index_sum_1_req_0;
      array_obj_ref_71_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_71_index_sum_1_req_1;
      array_obj_ref_71_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : array_obj_ref_56_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_56_load_0_req_0;
      array_obj_ref_56_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_56_load_0_req_1;
      array_obj_ref_56_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_56_word_address_0;
      array_obj_ref_56_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(7 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : array_obj_ref_61_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_61_load_0_req_0;
      array_obj_ref_61_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_61_load_0_req_1;
      array_obj_ref_61_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_61_word_address_0;
      array_obj_ref_61_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(7 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : array_obj_ref_66_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_66_load_0_req_0;
      array_obj_ref_66_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_66_load_0_req_1;
      array_obj_ref_66_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_66_word_address_0;
      array_obj_ref_66_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(7 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : array_obj_ref_71_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_71_load_0_req_0;
      array_obj_ref_71_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_71_load_0_req_1;
      array_obj_ref_71_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_71_word_address_0;
      array_obj_ref_71_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(7 downto 0),
          mtag => memory_space_3_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : array_obj_ref_75_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_75_load_0_req_0;
      array_obj_ref_75_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_75_load_0_req_1;
      array_obj_ref_75_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_75_word_address_0;
      array_obj_ref_75_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(2 downto 0),
          mtag => memory_space_4_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : array_obj_ref_79_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_79_load_0_req_0;
      array_obj_ref_79_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_79_load_0_req_1;
      array_obj_ref_79_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_79_word_address_0;
      array_obj_ref_79_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(2 downto 0),
          mtag => memory_space_5_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : array_obj_ref_83_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_83_load_0_req_0;
      array_obj_ref_83_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_83_load_0_req_1;
      array_obj_ref_83_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_83_word_address_0;
      array_obj_ref_83_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(2 downto 0),
          mtag => memory_space_6_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : array_obj_ref_87_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_87_load_0_req_0;
      array_obj_ref_87_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_87_load_0_req_1;
      array_obj_ref_87_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup7_gI: SplitGuardInterface generic map(name => "LoadGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_87_word_address_0;
      array_obj_ref_87_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup7", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(2 downto 0),
          mtag => memory_space_7_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup7 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(31 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- 
  end Block; -- data_path
  -- 
end dotP_even_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity dotP_odd is -- 
  generic (tag_length : integer); 
  port ( -- 
    R : in  std_logic_vector(7 downto 0);
    result : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity dotP_odd;
architecture dotP_odd_arch of dotP_odd is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal R_buffer :  std_logic_vector(7 downto 0);
  signal R_update_enable: Boolean;
  -- output port buffer signals
  signal result_buffer :  std_logic_vector(31 downto 0);
  signal result_update_enable: Boolean;
  signal dotP_odd_CP_995_start: Boolean;
  signal dotP_odd_CP_995_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nC_306_180_buf_req_1 : boolean;
  signal nval_1_266_190_buf_req_1 : boolean;
  signal ADD_u32_u32_319_inst_req_0 : boolean;
  signal nval_0_251_185_buf_ack_0 : boolean;
  signal phi_stmt_181_ack_0 : boolean;
  signal array_obj_ref_236_load_0_ack_0 : boolean;
  signal nC_306_180_buf_ack_1 : boolean;
  signal do_while_stmt_174_branch_ack_1 : boolean;
  signal W_val_3_267_delayed_5_0_287_inst_ack_1 : boolean;
  signal W_val_3_267_delayed_5_0_287_inst_req_1 : boolean;
  signal array_obj_ref_232_load_0_ack_1 : boolean;
  signal nC_306_180_buf_req_0 : boolean;
  signal ADD_u32_u32_319_inst_ack_0 : boolean;
  signal nC_306_180_buf_ack_0 : boolean;
  signal phi_stmt_186_req_1 : boolean;
  signal phi_stmt_181_req_1 : boolean;
  signal ADD_u8_u8_305_inst_req_1 : boolean;
  signal array_obj_ref_236_load_0_req_1 : boolean;
  signal array_obj_ref_232_load_0_ack_0 : boolean;
  signal array_obj_ref_232_load_0_req_0 : boolean;
  signal do_while_stmt_174_branch_ack_0 : boolean;
  signal ADD_u8_u8_305_inst_req_0 : boolean;
  signal array_obj_ref_236_load_0_req_0 : boolean;
  signal nval_0_251_185_buf_req_1 : boolean;
  signal nval_0_251_185_buf_ack_1 : boolean;
  signal array_obj_ref_232_load_0_req_1 : boolean;
  signal do_while_stmt_174_branch_req_0 : boolean;
  signal phi_stmt_176_ack_0 : boolean;
  signal array_obj_ref_236_load_0_ack_1 : boolean;
  signal phi_stmt_176_req_1 : boolean;
  signal ADD_u8_u8_305_inst_ack_1 : boolean;
  signal phi_stmt_181_req_0 : boolean;
  signal phi_stmt_176_req_0 : boolean;
  signal ADD_u32_u32_319_inst_req_1 : boolean;
  signal nval_1_266_190_buf_req_0 : boolean;
  signal nval_1_266_190_buf_ack_0 : boolean;
  signal ADD_u32_u32_319_inst_ack_1 : boolean;
  signal phi_stmt_191_req_1 : boolean;
  signal nval_1_266_190_buf_ack_1 : boolean;
  signal ADD_u8_u8_305_inst_ack_0 : boolean;
  signal phi_stmt_191_req_0 : boolean;
  signal W_val_3_267_delayed_5_0_287_inst_ack_0 : boolean;
  signal phi_stmt_186_ack_0 : boolean;
  signal W_val_2_255_delayed_5_0_272_inst_req_1 : boolean;
  signal phi_stmt_191_ack_0 : boolean;
  signal W_val_3_267_delayed_5_0_287_inst_req_0 : boolean;
  signal W_val_2_255_delayed_5_0_272_inst_ack_1 : boolean;
  signal W_val_1_243_delayed_5_0_257_inst_ack_1 : boolean;
  signal W_val_1_243_delayed_5_0_257_inst_req_1 : boolean;
  signal W_val_1_243_delayed_5_0_257_inst_ack_0 : boolean;
  signal nval_2_281_195_buf_req_0 : boolean;
  signal nval_2_281_195_buf_ack_0 : boolean;
  signal nval_2_281_195_buf_req_1 : boolean;
  signal nval_2_281_195_buf_ack_1 : boolean;
  signal array_obj_ref_228_load_0_ack_1 : boolean;
  signal W_val_1_243_delayed_5_0_257_inst_req_0 : boolean;
  signal W_val_2_255_delayed_5_0_272_inst_req_0 : boolean;
  signal W_val_2_255_delayed_5_0_272_inst_ack_0 : boolean;
  signal phi_stmt_186_req_0 : boolean;
  signal nval_0_251_185_buf_req_0 : boolean;
  signal W_val_0_231_delayed_5_0_242_inst_ack_1 : boolean;
  signal W_val_0_231_delayed_5_0_242_inst_req_1 : boolean;
  signal phi_stmt_196_req_1 : boolean;
  signal phi_stmt_196_req_0 : boolean;
  signal W_val_0_231_delayed_5_0_242_inst_ack_0 : boolean;
  signal W_val_0_231_delayed_5_0_242_inst_req_0 : boolean;
  signal phi_stmt_196_ack_0 : boolean;
  signal array_obj_ref_240_load_0_ack_1 : boolean;
  signal array_obj_ref_240_load_0_req_1 : boolean;
  signal array_obj_ref_240_load_0_ack_0 : boolean;
  signal array_obj_ref_240_load_0_req_0 : boolean;
  signal nval_3_296_200_buf_req_0 : boolean;
  signal nval_3_296_200_buf_ack_0 : boolean;
  signal nval_3_296_200_buf_req_1 : boolean;
  signal nval_3_296_200_buf_ack_1 : boolean;
  signal array_obj_ref_228_load_0_req_1 : boolean;
  signal array_obj_ref_209_index_0_scale_req_0 : boolean;
  signal array_obj_ref_209_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_209_index_0_scale_req_1 : boolean;
  signal array_obj_ref_209_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_209_index_sum_1_req_0 : boolean;
  signal array_obj_ref_209_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_209_index_sum_1_req_1 : boolean;
  signal array_obj_ref_209_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_209_load_0_req_0 : boolean;
  signal array_obj_ref_209_load_0_ack_0 : boolean;
  signal array_obj_ref_209_load_0_req_1 : boolean;
  signal array_obj_ref_209_load_0_ack_1 : boolean;
  signal array_obj_ref_214_index_0_scale_req_0 : boolean;
  signal array_obj_ref_214_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_214_index_0_scale_req_1 : boolean;
  signal array_obj_ref_214_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_214_index_sum_1_req_0 : boolean;
  signal array_obj_ref_214_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_214_index_sum_1_req_1 : boolean;
  signal array_obj_ref_214_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_214_load_0_req_0 : boolean;
  signal array_obj_ref_214_load_0_ack_0 : boolean;
  signal array_obj_ref_214_load_0_req_1 : boolean;
  signal array_obj_ref_214_load_0_ack_1 : boolean;
  signal array_obj_ref_219_index_0_scale_req_0 : boolean;
  signal array_obj_ref_219_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_219_index_0_scale_req_1 : boolean;
  signal array_obj_ref_219_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_219_index_sum_1_req_0 : boolean;
  signal array_obj_ref_219_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_219_index_sum_1_req_1 : boolean;
  signal array_obj_ref_219_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_219_load_0_req_0 : boolean;
  signal array_obj_ref_219_load_0_ack_0 : boolean;
  signal array_obj_ref_219_load_0_req_1 : boolean;
  signal array_obj_ref_219_load_0_ack_1 : boolean;
  signal array_obj_ref_224_index_0_scale_req_0 : boolean;
  signal array_obj_ref_224_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_224_index_0_scale_req_1 : boolean;
  signal array_obj_ref_224_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_224_index_sum_1_req_0 : boolean;
  signal array_obj_ref_224_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_224_index_sum_1_req_1 : boolean;
  signal array_obj_ref_224_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_224_load_0_req_0 : boolean;
  signal array_obj_ref_224_load_0_ack_0 : boolean;
  signal array_obj_ref_224_load_0_req_1 : boolean;
  signal array_obj_ref_224_load_0_ack_1 : boolean;
  signal array_obj_ref_228_load_0_req_0 : boolean;
  signal array_obj_ref_228_load_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "dotP_odd_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 8) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= R;
  R_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(tag_length + 7 downto 8) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 7 downto 8);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  dotP_odd_CP_995_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "dotP_odd_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= result_buffer;
  result <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= dotP_odd_CP_995_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= dotP_odd_CP_995_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= dotP_odd_CP_995_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  dotP_odd_CP_995: Block -- control-path 
    signal dotP_odd_CP_995_elements: BooleanArray(202 downto 0);
    -- 
  begin -- 
    dotP_odd_CP_995_elements(0) <= dotP_odd_CP_995_start;
    dotP_odd_CP_995_symbol <= dotP_odd_CP_995_elements(202);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_173/$entry
      -- CP-element group 0: 	 branch_block_stmt_173/branch_block_stmt_173__entry__
      -- CP-element group 0: 	 branch_block_stmt_173/do_while_stmt_174__entry__
      -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	200 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	202 
    -- CP-element group 1: 	201 
    -- CP-element group 1:  members (10) 
      -- CP-element group 1: 	 assign_stmt_320/$entry
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_Sample/rr
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_update_start_
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_173/$exit
      -- CP-element group 1: 	 branch_block_stmt_173/branch_block_stmt_173__exit__
      -- CP-element group 1: 	 branch_block_stmt_173/do_while_stmt_174__exit__
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_Update/cr
      -- CP-element group 1: 	 assign_stmt_320/ADD_u32_u32_319_Update/$entry
      -- 
    rr_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(1), ack => ADD_u32_u32_319_inst_req_0); -- 
    cr_1988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(1), ack => ADD_u32_u32_319_inst_req_1); -- 
    dotP_odd_CP_995_elements(1) <= dotP_odd_CP_995_elements(200);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_173/do_while_stmt_174/$entry
      -- CP-element group 2: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174__entry__
      -- 
    dotP_odd_CP_995_elements(2) <= dotP_odd_CP_995_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	200 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174__exit__
      -- 
    -- Element group dotP_odd_CP_995_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_173/do_while_stmt_174/loop_back
      -- 
    -- Element group dotP_odd_CP_995_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	198 
    -- CP-element group 5: 	199 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_173/do_while_stmt_174/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_173/do_while_stmt_174/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_173/do_while_stmt_174/condition_done
      -- 
    dotP_odd_CP_995_elements(5) <= dotP_odd_CP_995_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	197 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_173/do_while_stmt_174/loop_body_done
      -- 
    dotP_odd_CP_995_elements(6) <= dotP_odd_CP_995_elements(197);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	95 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/back_edge_to_loop_body
      -- 
    dotP_odd_CP_995_elements(7) <= dotP_odd_CP_995_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	97 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/first_time_through_loop_body
      -- 
    dotP_odd_CP_995_elements(8) <= dotP_odd_CP_995_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	142 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	196 
    -- CP-element group 9: 	151 
    -- CP-element group 9: 	125 
    -- CP-element group 9: 	124 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	90 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	112 
    -- CP-element group 9: 	116 
    -- CP-element group 9:  members (26) 
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_0/index_resize_ack
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resized_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_computed_0
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_0/index_resize_req
      -- CP-element group 9: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_0/index_resize_ack
      -- 
    -- Element group dotP_odd_CP_995_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	195 
    -- CP-element group 10: 	196 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/condition_evaluated
      -- 
    condition_evaluated_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(10), ack => do_while_stmt_174_branch_req_0); -- 
    dotP_odd_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(14) & dotP_odd_CP_995_elements(195) & dotP_odd_CP_995_elements(196);
      gj_dotP_odd_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	89 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	91 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_sample_start__ps
      -- 
    dotP_odd_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(15) & dotP_odd_CP_995_elements(32) & dotP_odd_CP_995_elements(51) & dotP_odd_CP_995_elements(70) & dotP_odd_CP_995_elements(89) & dotP_odd_CP_995_elements(14);
      gj_dotP_odd_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	92 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	148 
    -- CP-element group 12: 	177 
    -- CP-element group 12: 	181 
    -- CP-element group 12: 	169 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	173 
    -- CP-element group 12: 	122 
    -- CP-element group 12: 	185 
    -- CP-element group 12: 	189 
    -- CP-element group 12: 	193 
    -- CP-element group 12: 	161 
    -- CP-element group 12: 	165 
    -- CP-element group 12: 	109 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	89 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_sample_completed_
      -- 
    dotP_odd_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(17) & dotP_odd_CP_995_elements(35) & dotP_odd_CP_995_elements(54) & dotP_odd_CP_995_elements(73) & dotP_odd_CP_995_elements(92);
      gj_dotP_odd_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	90 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	93 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/aggregated_phi_update_req
      -- 
    dotP_odd_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(16) & dotP_odd_CP_995_elements(33) & dotP_odd_CP_995_elements(52) & dotP_odd_CP_995_elements(71) & dotP_odd_CP_995_elements(90);
      gj_dotP_odd_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	94 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/aggregated_phi_update_ack
      -- 
    dotP_odd_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(37) & dotP_odd_CP_995_elements(56) & dotP_odd_CP_995_elements(75) & dotP_odd_CP_995_elements(94);
      gj_dotP_odd_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: 	195 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_sample_start_
      -- 
    dotP_odd_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(195);
      gj_dotP_odd_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	162 
    -- CP-element group 16: 	170 
    -- CP-element group 16: 	166 
    -- CP-element group 16: 	156 
    -- CP-element group 16: 	143 
    -- CP-element group 16: 	130 
    -- CP-element group 16: 	174 
    -- CP-element group 16: 	194 
    -- CP-element group 16: 	117 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_update_start_
      -- 
    dotP_odd_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1,7 => 0,8 => 0,9 => 1);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(162) & dotP_odd_CP_995_elements(170) & dotP_odd_CP_995_elements(166) & dotP_odd_CP_995_elements(156) & dotP_odd_CP_995_elements(143) & dotP_odd_CP_995_elements(130) & dotP_odd_CP_995_elements(174) & dotP_odd_CP_995_elements(194) & dotP_odd_CP_995_elements(117);
      gj_dotP_odd_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_sample_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	164 
    -- CP-element group 18: 	168 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	154 
    -- CP-element group 18: 	141 
    -- CP-element group 18: 	172 
    -- CP-element group 18: 	128 
    -- CP-element group 18: 	192 
    -- CP-element group 18: 	160 
    -- CP-element group 18: 	115 
    -- CP-element group 18:  members (150) 
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_word_addrgen/root_register_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resized_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scaled_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_computed_1
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_1/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_resize_1/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_1/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_1/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_1/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_1/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_word_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_resized_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_scaled_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_computed_0
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_resize_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_resize_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_resize_0/index_resize_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_resize_0/index_resize_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_scale_0/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_scale_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_scale_0/scale_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_index_scale_0/scale_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_final_index_sum_regn/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_final_index_sum_regn/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_final_index_sum_regn/req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_final_index_sum_regn/ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_word_addrgen/$entry
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_word_addrgen/$exit
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_word_addrgen/root_register_req
      -- CP-element group 18: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_word_addrgen/root_register_ack
      -- 
    -- Element group dotP_odd_CP_995_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_loopback_trigger
      -- 
    dotP_odd_CP_995_elements(19) <= dotP_odd_CP_995_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_loopback_sample_req
      -- 
    phi_stmt_176_loopback_sample_req_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_176_loopback_sample_req_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(20), ack => phi_stmt_176_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_entry_trigger
      -- 
    dotP_odd_CP_995_elements(21) <= dotP_odd_CP_995_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_entry_sample_req
      -- 
    phi_stmt_176_entry_sample_req_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_176_entry_sample_req_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(22), ack => phi_stmt_176_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_176_phi_mux_ack_ps
      -- 
    phi_stmt_176_phi_mux_ack_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_176_ack_0, ack => dotP_odd_CP_995_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_sample_start__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_update_start_
      -- CP-element group 25: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_update_start__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_update_completed__ps
      -- 
    dotP_odd_CP_995_elements(26) <= dotP_odd_CP_995_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_179_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(25), ack => dotP_odd_CP_995_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_sample_start_
      -- 
    req_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(28), ack => nC_306_180_buf_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Update/req
      -- CP-element group 29: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_update_start_
      -- CP-element group 29: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Update/$entry
      -- 
    req_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(29), ack => nC_306_180_buf_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_sample_completed_
      -- 
    ack_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nC_306_180_buf_ack_0, ack => dotP_odd_CP_995_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nC_180_Update/$exit
      -- 
    ack_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nC_306_180_buf_ack_1, ack => dotP_odd_CP_995_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	163 
    -- CP-element group 32: 	12 
    -- CP-element group 32: 	179 
    -- CP-element group 32: 	120 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_sample_start_
      -- 
    dotP_odd_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(163) & dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(179) & dotP_odd_CP_995_elements(120);
      gj_dotP_odd_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	178 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_update_start_
      -- 
    dotP_odd_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(178);
      gj_dotP_odd_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_sample_start__ps
      -- 
    dotP_odd_CP_995_elements(34) <= dotP_odd_CP_995_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_sample_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_update_start__ps
      -- 
    dotP_odd_CP_995_elements(36) <= dotP_odd_CP_995_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	176 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_loopback_trigger
      -- 
    dotP_odd_CP_995_elements(38) <= dotP_odd_CP_995_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_loopback_sample_req_ps
      -- 
    phi_stmt_181_loopback_sample_req_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_181_loopback_sample_req_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(39), ack => phi_stmt_181_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_entry_trigger
      -- 
    dotP_odd_CP_995_elements(40) <= dotP_odd_CP_995_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_entry_sample_req_ps
      -- 
    phi_stmt_181_entry_sample_req_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_181_entry_sample_req_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(41), ack => phi_stmt_181_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_181_phi_mux_ack_ps
      -- 
    phi_stmt_181_phi_mux_ack_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_181_ack_0, ack => dotP_odd_CP_995_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_sample_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_update_start_
      -- 
    -- Element group dotP_odd_CP_995_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_update_completed__ps
      -- 
    dotP_odd_CP_995_elements(45) <= dotP_odd_CP_995_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_184_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(44), ack => dotP_odd_CP_995_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Sample/req
      -- 
    req_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(47), ack => nval_0_251_185_buf_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_update_start_
      -- CP-element group 48: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Update/req
      -- 
    req_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(48), ack => nval_0_251_185_buf_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Sample/$exit
      -- 
    ack_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_0_251_185_buf_ack_0, ack => dotP_odd_CP_995_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_0_185_Update/ack
      -- 
    ack_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_0_251_185_buf_ack_1, ack => dotP_odd_CP_995_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	167 
    -- CP-element group 51: 	12 
    -- CP-element group 51: 	183 
    -- CP-element group 51: 	133 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_sample_start_
      -- 
    dotP_odd_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(167) & dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(183) & dotP_odd_CP_995_elements(133);
      gj_dotP_odd_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	182 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_update_start_
      -- 
    dotP_odd_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(182);
      gj_dotP_odd_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_sample_start__ps
      -- 
    dotP_odd_CP_995_elements(53) <= dotP_odd_CP_995_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_sample_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_update_start__ps
      -- 
    dotP_odd_CP_995_elements(55) <= dotP_odd_CP_995_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	180 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_loopback_trigger
      -- 
    dotP_odd_CP_995_elements(57) <= dotP_odd_CP_995_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_loopback_sample_req_ps
      -- 
    phi_stmt_186_loopback_sample_req_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_186_loopback_sample_req_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(58), ack => phi_stmt_186_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_entry_trigger
      -- 
    dotP_odd_CP_995_elements(59) <= dotP_odd_CP_995_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_entry_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_entry_sample_req
      -- 
    phi_stmt_186_entry_sample_req_1125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_186_entry_sample_req_1125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(60), ack => phi_stmt_186_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_phi_mux_ack_ps
      -- CP-element group 61: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_186_phi_mux_ack
      -- 
    phi_stmt_186_phi_mux_ack_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_186_ack_0, ack => dotP_odd_CP_995_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_sample_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_update_start_
      -- 
    -- Element group dotP_odd_CP_995_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_update_completed__ps
      -- 
    dotP_odd_CP_995_elements(64) <= dotP_odd_CP_995_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_189_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(63), ack => dotP_odd_CP_995_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Sample/$entry
      -- 
    req_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(66), ack => nval_1_266_190_buf_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Update/req
      -- CP-element group 67: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_update_start_
      -- CP-element group 67: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Update/$entry
      -- 
    req_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(67), ack => nval_1_266_190_buf_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_sample_completed_
      -- 
    ack_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_1_266_190_buf_ack_0, ack => dotP_odd_CP_995_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_1_190_Update/ack
      -- 
    ack_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_1_266_190_buf_ack_1, ack => dotP_odd_CP_995_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	171 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	146 
    -- CP-element group 70: 	187 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_sample_start_
      -- 
    dotP_odd_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(171) & dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(146) & dotP_odd_CP_995_elements(187);
      gj_dotP_odd_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	186 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_update_start_
      -- 
    dotP_odd_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(186);
      gj_dotP_odd_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_sample_start__ps
      -- 
    dotP_odd_CP_995_elements(72) <= dotP_odd_CP_995_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_sample_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_update_start__ps
      -- 
    dotP_odd_CP_995_elements(74) <= dotP_odd_CP_995_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	184 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_loopback_trigger
      -- 
    dotP_odd_CP_995_elements(76) <= dotP_odd_CP_995_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_loopback_sample_req_ps
      -- CP-element group 77: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_loopback_sample_req
      -- 
    phi_stmt_191_loopback_sample_req_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_191_loopback_sample_req_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(77), ack => phi_stmt_191_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_entry_trigger
      -- 
    dotP_odd_CP_995_elements(78) <= dotP_odd_CP_995_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_entry_sample_req_ps
      -- 
    phi_stmt_191_entry_sample_req_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_191_entry_sample_req_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(79), ack => phi_stmt_191_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_191_phi_mux_ack
      -- 
    phi_stmt_191_phi_mux_ack_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_191_ack_0, ack => dotP_odd_CP_995_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_sample_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_update_start_
      -- 
    -- Element group dotP_odd_CP_995_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_update_completed__ps
      -- 
    dotP_odd_CP_995_elements(83) <= dotP_odd_CP_995_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_194_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(82), ack => dotP_odd_CP_995_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Sample/req
      -- 
    req_1193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(85), ack => nval_2_281_195_buf_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_update_start_
      -- CP-element group 86: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Update/req
      -- 
    req_1198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(86), ack => nval_2_281_195_buf_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Sample/ack
      -- 
    ack_1194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_2_281_195_buf_ack_0, ack => dotP_odd_CP_995_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_2_195_Update/ack
      -- 
    ack_1199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_2_281_195_buf_ack_1, ack => dotP_odd_CP_995_elements(88)); -- 
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	12 
    -- CP-element group 89: 	175 
    -- CP-element group 89: 	191 
    -- CP-element group 89: 	159 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	11 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_sample_start_
      -- 
    dotP_odd_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(175) & dotP_odd_CP_995_elements(191) & dotP_odd_CP_995_elements(159);
      gj_dotP_odd_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	9 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	190 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	13 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_update_start_
      -- 
    dotP_odd_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "dotP_odd_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(190);
      gj_dotP_odd_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	11 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_sample_start__ps
      -- 
    dotP_odd_CP_995_elements(91) <= dotP_odd_CP_995_elements(11);
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	12 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_sample_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(92) is bound as output of CP function.
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	13 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_update_start__ps
      -- 
    dotP_odd_CP_995_elements(93) <= dotP_odd_CP_995_elements(13);
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: 	188 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_update_completed__ps
      -- 
    -- Element group dotP_odd_CP_995_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	7 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_loopback_trigger
      -- 
    dotP_odd_CP_995_elements(95) <= dotP_odd_CP_995_elements(7);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_loopback_sample_req
      -- CP-element group 96: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_loopback_sample_req_ps
      -- 
    phi_stmt_196_loopback_sample_req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_196_loopback_sample_req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(96), ack => phi_stmt_196_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	8 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_entry_trigger
      -- 
    dotP_odd_CP_995_elements(97) <= dotP_odd_CP_995_elements(8);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_entry_sample_req
      -- CP-element group 98: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_entry_sample_req_ps
      -- 
    phi_stmt_196_entry_sample_req_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_196_entry_sample_req_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(98), ack => phi_stmt_196_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_phi_mux_ack
      -- CP-element group 99: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/phi_stmt_196_phi_mux_ack_ps
      -- 
    phi_stmt_196_phi_mux_ack_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_196_ack_0, ack => dotP_odd_CP_995_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_sample_completed__ps
      -- CP-element group 100: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_sample_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_update_start_
      -- 
    -- Element group dotP_odd_CP_995_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_update_completed__ps
      -- 
    dotP_odd_CP_995_elements(102) <= dotP_odd_CP_995_elements(103);
    -- CP-element group 103:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	102 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/type_cast_199_update_completed_
      -- 
    -- Element group dotP_odd_CP_995_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(101), ack => dotP_odd_CP_995_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Sample/req
      -- 
    req_1237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(104), ack => nval_3_296_200_buf_req_0); -- 
    -- Element group dotP_odd_CP_995_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_update_start_
      -- CP-element group 105: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Update/req
      -- 
    req_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(105), ack => nval_3_296_200_buf_req_1); -- 
    -- Element group dotP_odd_CP_995_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Sample/ack
      -- 
    ack_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_3_296_200_buf_ack_0, ack => dotP_odd_CP_995_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/R_nval_3_200_Update/ack
      -- 
    ack_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nval_3_296_200_buf_ack_1, ack => dotP_odd_CP_995_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	118 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	119 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/word_0/rr
      -- 
    rr_1326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(108), ack => array_obj_ref_209_load_0_req_0); -- 
    dotP_odd_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(118) & dotP_odd_CP_995_elements(119);
      gj_dotP_odd_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	12 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	120 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	120 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_update_start_
      -- CP-element group 109: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/$entry
      -- CP-element group 109: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/word_0/cr
      -- 
    cr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(109), ack => array_obj_ref_209_load_0_req_1); -- 
    dotP_odd_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(120);
      gj_dotP_odd_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	114 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	117 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	115 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scaled_0
      -- 
    dotP_odd_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(114) & dotP_odd_CP_995_elements(117);
      gj_dotP_odd_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_sample_start
      -- CP-element group 111: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Sample/rr
      -- 
    rr_1268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(111), ack => array_obj_ref_209_index_0_scale_req_0); -- 
    dotP_odd_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(113);
      gj_dotP_odd_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	9 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_update_start
      -- CP-element group 112: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Update/cr
      -- 
    cr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(112), ack => array_obj_ref_209_index_0_scale_req_1); -- 
    dotP_odd_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(114);
      gj_dotP_odd_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	197 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_sample_complete
      -- CP-element group 113: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Sample/ra
      -- 
    ra_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_index_0_scale_ack_0, ack => dotP_odd_CP_995_elements(113)); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	110 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_update_complete
      -- CP-element group 114: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_index_scale_0_Update/ca
      -- 
    ca_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_index_0_scale_ack_1, ack => dotP_odd_CP_995_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	18 
    -- CP-element group 115: 	110 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_sample_start
      -- CP-element group 115: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Sample/rr
      -- 
    rr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(115), ack => array_obj_ref_209_index_sum_1_req_0); -- 
    dotP_odd_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(110) & dotP_odd_CP_995_elements(117);
      gj_dotP_odd_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	119 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_update_start
      -- CP-element group 116: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Update/cr
      -- 
    cr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(116), ack => array_obj_ref_209_index_sum_1_req_1); -- 
    dotP_odd_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(119);
      gj_dotP_odd_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	197 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	16 
    -- CP-element group 117: 	110 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_sample_complete
      -- CP-element group 117: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Sample/ra
      -- 
    ra_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_index_sum_1_ack_0, ack => dotP_odd_CP_995_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	108 
    -- CP-element group 118:  members (18) 
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_word_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_root_address_calculated
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_offset_calculated
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_update_complete
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_partial_sum_1_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_final_index_sum_regn/$entry
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_final_index_sum_regn/$exit
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_final_index_sum_regn/req
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_final_index_sum_regn/ack
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_base_plus_offset/$entry
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_base_plus_offset/$exit
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_base_plus_offset/sum_rename_req
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_base_plus_offset/sum_rename_ack
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_word_addrgen/$entry
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_word_addrgen/$exit
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_word_addrgen/root_register_req
      -- CP-element group 118: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_word_addrgen/root_register_ack
      -- 
    ca_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_index_sum_1_ack_1, ack => dotP_odd_CP_995_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	116 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Sample/word_access_start/word_0/ra
      -- 
    ra_1327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_load_0_ack_0, ack => dotP_odd_CP_995_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	109 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	197 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	32 
    -- CP-element group 120: 	109 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/array_obj_ref_209_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/array_obj_ref_209_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/array_obj_ref_209_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_209_Update/array_obj_ref_209_Merge/merge_ack
      -- 
    ca_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_209_load_0_ack_1, ack => dotP_odd_CP_995_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	131 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	132 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	132 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/$entry
      -- CP-element group 121: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/word_0/$entry
      -- CP-element group 121: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/word_0/rr
      -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(121), ack => array_obj_ref_214_load_0_req_0); -- 
    dotP_odd_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(131) & dotP_odd_CP_995_elements(132);
      gj_dotP_odd_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	12 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	133 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	133 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_update_start_
      -- CP-element group 122: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/$entry
      -- CP-element group 122: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/word_0/$entry
      -- CP-element group 122: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/word_0/cr
      -- 
    cr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(122), ack => array_obj_ref_214_load_0_req_1); -- 
    dotP_odd_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(133);
      gj_dotP_odd_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	130 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scaled_0
      -- 
    dotP_odd_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(127) & dotP_odd_CP_995_elements(130);
      gj_dotP_odd_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	9 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_sample_start
      -- CP-element group 124: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Sample/rr
      -- 
    rr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(124), ack => array_obj_ref_214_index_0_scale_req_0); -- 
    dotP_odd_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(126);
      gj_dotP_odd_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	9 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_update_start
      -- CP-element group 125: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Update/cr
      -- 
    cr_1372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(125), ack => array_obj_ref_214_index_0_scale_req_1); -- 
    dotP_odd_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(127);
      gj_dotP_odd_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	197 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Sample/ra
      -- 
    ra_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_index_0_scale_ack_0, ack => dotP_odd_CP_995_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_update_complete
      -- CP-element group 127: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_index_scale_0_Update/ca
      -- 
    ca_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_index_0_scale_ack_1, ack => dotP_odd_CP_995_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	18 
    -- CP-element group 128: 	123 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_sample_start
      -- CP-element group 128: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Sample/rr
      -- 
    rr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(128), ack => array_obj_ref_214_index_sum_1_req_0); -- 
    dotP_odd_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(123) & dotP_odd_CP_995_elements(130);
      gj_dotP_odd_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	132 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_update_start
      -- CP-element group 129: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Update/cr
      -- 
    cr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(129), ack => array_obj_ref_214_index_sum_1_req_1); -- 
    dotP_odd_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(132);
      gj_dotP_odd_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	197 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	16 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	123 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_sample_complete
      -- CP-element group 130: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Sample/ra
      -- 
    ra_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_index_sum_1_ack_0, ack => dotP_odd_CP_995_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	121 
    -- CP-element group 131:  members (18) 
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_word_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_root_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_offset_calculated
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_update_complete
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_partial_sum_1_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_final_index_sum_regn/$entry
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_final_index_sum_regn/$exit
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_final_index_sum_regn/req
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_final_index_sum_regn/ack
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_base_plus_offset/$entry
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_base_plus_offset/$exit
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_base_plus_offset/sum_rename_req
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_base_plus_offset/sum_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_word_addrgen/$entry
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_word_addrgen/$exit
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_word_addrgen/root_register_req
      -- CP-element group 131: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_word_addrgen/root_register_ack
      -- 
    ca_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_index_sum_1_ack_1, ack => dotP_odd_CP_995_elements(131)); -- 
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	121 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	129 
    -- CP-element group 132: 	121 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/$exit
      -- CP-element group 132: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/word_0/$exit
      -- CP-element group 132: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Sample/word_access_start/word_0/ra
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_load_0_ack_0, ack => dotP_odd_CP_995_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	122 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	197 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	122 
    -- CP-element group 133: 	51 
    -- CP-element group 133:  members (9) 
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/$exit
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/word_0/$exit
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/word_access_complete/word_0/ca
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/array_obj_ref_214_Merge/$entry
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/array_obj_ref_214_Merge/$exit
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/array_obj_ref_214_Merge/merge_req
      -- CP-element group 133: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_214_Update/array_obj_ref_214_Merge/merge_ack
      -- 
    ca_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_214_load_0_ack_1, ack => dotP_odd_CP_995_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	144 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	145 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	145 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/$entry
      -- CP-element group 134: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/word_0/rr
      -- 
    rr_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(134), ack => array_obj_ref_219_load_0_req_0); -- 
    dotP_odd_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(144) & dotP_odd_CP_995_elements(145);
      gj_dotP_odd_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	146 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	146 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_update_start_
      -- CP-element group 135: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/$entry
      -- CP-element group 135: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/word_0/$entry
      -- CP-element group 135: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/word_0/cr
      -- 
    cr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(135), ack => array_obj_ref_219_load_0_req_1); -- 
    dotP_odd_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(146);
      gj_dotP_odd_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	140 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	143 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scaled_0
      -- 
    dotP_odd_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(140) & dotP_odd_CP_995_elements(143);
      gj_dotP_odd_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_sample_start
      -- CP-element group 137: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Sample/rr
      -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(137), ack => array_obj_ref_219_index_0_scale_req_0); -- 
    dotP_odd_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(139);
      gj_dotP_odd_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_update_start
      -- CP-element group 138: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Update/cr
      -- 
    cr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(138), ack => array_obj_ref_219_index_0_scale_req_1); -- 
    dotP_odd_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(140);
      gj_dotP_odd_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	197 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_sample_complete
      -- CP-element group 139: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Sample/ra
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_index_0_scale_ack_0, ack => dotP_odd_CP_995_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	136 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_update_complete
      -- CP-element group 140: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_index_scale_0_Update/ca
      -- 
    ca_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_index_0_scale_ack_1, ack => dotP_odd_CP_995_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	18 
    -- CP-element group 141: 	136 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_sample_start
      -- CP-element group 141: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Sample/rr
      -- 
    rr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(141), ack => array_obj_ref_219_index_sum_1_req_0); -- 
    dotP_odd_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(136) & dotP_odd_CP_995_elements(143);
      gj_dotP_odd_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	9 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	145 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_update_start
      -- CP-element group 142: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Update/cr
      -- 
    cr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(142), ack => array_obj_ref_219_index_sum_1_req_1); -- 
    dotP_odd_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(145);
      gj_dotP_odd_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	197 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	16 
    -- CP-element group 143: 	141 
    -- CP-element group 143: 	136 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_sample_complete
      -- CP-element group 143: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Sample/ra
      -- 
    ra_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_index_sum_1_ack_0, ack => dotP_odd_CP_995_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	134 
    -- CP-element group 144:  members (18) 
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_root_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_offset_calculated
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_word_address_calculated
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_update_complete
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_partial_sum_1_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_final_index_sum_regn/$entry
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_final_index_sum_regn/$exit
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_final_index_sum_regn/req
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_final_index_sum_regn/ack
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_base_plus_offset/$entry
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_base_plus_offset/$exit
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_base_plus_offset/sum_rename_req
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_base_plus_offset/sum_rename_ack
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_word_addrgen/$entry
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_word_addrgen/$exit
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_word_addrgen/root_register_req
      -- CP-element group 144: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_word_addrgen/root_register_ack
      -- 
    ca_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_index_sum_1_ack_1, ack => dotP_odd_CP_995_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	134 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: 	134 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Sample/word_access_start/word_0/ra
      -- 
    ra_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_load_0_ack_0, ack => dotP_odd_CP_995_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	135 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	197 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	135 
    -- CP-element group 146: 	70 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/array_obj_ref_219_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/array_obj_ref_219_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/array_obj_ref_219_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_219_Update/array_obj_ref_219_Merge/merge_ack
      -- 
    ca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_219_load_0_ack_1, ack => dotP_odd_CP_995_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	157 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	158 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	158 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/$entry
      -- CP-element group 147: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/word_0/$entry
      -- CP-element group 147: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/word_0/rr
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(147), ack => array_obj_ref_224_load_0_req_0); -- 
    dotP_odd_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(157) & dotP_odd_CP_995_elements(158);
      gj_dotP_odd_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	12 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	159 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	159 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_update_start_
      -- CP-element group 148: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/$entry
      -- CP-element group 148: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/word_0/$entry
      -- CP-element group 148: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/word_0/cr
      -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(148), ack => array_obj_ref_224_load_0_req_1); -- 
    dotP_odd_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(159);
      gj_dotP_odd_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	153 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	156 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scaled_0
      -- 
    dotP_odd_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(153) & dotP_odd_CP_995_elements(156);
      gj_dotP_odd_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_sample_start
      -- CP-element group 150: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Sample/rr
      -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(150), ack => array_obj_ref_224_index_0_scale_req_0); -- 
    dotP_odd_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(152);
      gj_dotP_odd_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	9 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_update_start
      -- CP-element group 151: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Update/cr
      -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(151), ack => array_obj_ref_224_index_0_scale_req_1); -- 
    dotP_odd_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(153);
      gj_dotP_odd_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	197 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_sample_complete
      -- CP-element group 152: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Sample/ra
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_index_0_scale_ack_0, ack => dotP_odd_CP_995_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	149 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_update_complete
      -- CP-element group 153: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_index_scale_0_Update/ca
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_index_0_scale_ack_1, ack => dotP_odd_CP_995_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	18 
    -- CP-element group 154: 	149 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_sample_start
      -- CP-element group 154: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Sample/rr
      -- 
    rr_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(154), ack => array_obj_ref_224_index_sum_1_req_0); -- 
    dotP_odd_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(149) & dotP_odd_CP_995_elements(156);
      gj_dotP_odd_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	158 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_update_start
      -- CP-element group 155: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Update/cr
      -- 
    cr_1597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(155), ack => array_obj_ref_224_index_sum_1_req_1); -- 
    dotP_odd_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(9) & dotP_odd_CP_995_elements(158);
      gj_dotP_odd_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	197 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	16 
    -- CP-element group 156: 	154 
    -- CP-element group 156: 	149 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_sample_complete
      -- CP-element group 156: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Sample/ra
      -- 
    ra_1593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_index_sum_1_ack_0, ack => dotP_odd_CP_995_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	147 
    -- CP-element group 157:  members (18) 
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_word_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_root_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_offset_calculated
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_update_complete
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_partial_sum_1_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_final_index_sum_regn/$entry
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_final_index_sum_regn/$exit
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_final_index_sum_regn/req
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_final_index_sum_regn/ack
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_base_plus_offset/$entry
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_base_plus_offset/$exit
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_base_plus_offset/sum_rename_req
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_base_plus_offset/sum_rename_ack
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_word_addrgen/$entry
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_word_addrgen/$exit
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_word_addrgen/root_register_req
      -- CP-element group 157: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_word_addrgen/root_register_ack
      -- 
    ca_1598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_index_sum_1_ack_1, ack => dotP_odd_CP_995_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	147 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	147 
    -- CP-element group 158: 	155 
    -- CP-element group 158:  members (5) 
      -- CP-element group 158: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/$exit
      -- CP-element group 158: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Sample/word_access_start/word_0/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_load_0_ack_0, ack => dotP_odd_CP_995_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	148 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	197 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	148 
    -- CP-element group 159: 	89 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/$exit
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/word_0/$exit
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/word_access_complete/word_0/ca
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/array_obj_ref_224_Merge/$entry
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/array_obj_ref_224_Merge/$exit
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/array_obj_ref_224_Merge/merge_req
      -- CP-element group 159: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_224_Update/array_obj_ref_224_Merge/merge_ack
      -- 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_224_load_0_ack_1, ack => dotP_odd_CP_995_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	18 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/$entry
      -- CP-element group 160: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/word_0/rr
      -- 
    rr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(160), ack => array_obj_ref_228_load_0_req_0); -- 
    dotP_odd_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(162);
      gj_dotP_odd_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	12 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/word_0/cr
      -- CP-element group 161: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_update_start_
      -- CP-element group 161: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/$entry
      -- CP-element group 161: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/word_0/$entry
      -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(161), ack => array_obj_ref_228_load_0_req_1); -- 
    dotP_odd_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(163);
      gj_dotP_odd_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	16 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Sample/word_access_start/word_0/ra
      -- 
    ra_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_228_load_0_ack_0, ack => dotP_odd_CP_995_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	197 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	32 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/array_obj_ref_228_Merge/merge_ack
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/array_obj_ref_228_Merge/$exit
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/array_obj_ref_228_Merge/merge_req
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/array_obj_ref_228_Merge/$entry
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_228_Update/word_access_complete/$exit
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_228_load_0_ack_1, ack => dotP_odd_CP_995_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	18 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/word_0/$entry
      -- CP-element group 164: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/word_0/rr
      -- CP-element group 164: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/$entry
      -- 
    rr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(164), ack => array_obj_ref_232_load_0_req_0); -- 
    dotP_odd_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(166);
      gj_dotP_odd_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	12 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/$entry
      -- CP-element group 165: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/word_0/$entry
      -- CP-element group 165: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/word_0/cr
      -- CP-element group 165: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_update_start_
      -- CP-element group 165: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/$entry
      -- 
    cr_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(165), ack => array_obj_ref_232_load_0_req_1); -- 
    dotP_odd_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(167);
      gj_dotP_odd_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: 	16 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/word_0/$exit
      -- CP-element group 166: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/$exit
      -- CP-element group 166: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Sample/word_access_start/word_0/ra
      -- CP-element group 166: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_sample_completed_
      -- 
    ra_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_232_load_0_ack_0, ack => dotP_odd_CP_995_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	197 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: 	51 
    -- CP-element group 167:  members (9) 
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/array_obj_ref_232_Merge/$exit
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/$exit
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/array_obj_ref_232_Merge/$entry
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/word_0/ca
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/array_obj_ref_232_Merge/merge_ack
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/word_access_complete/word_0/$exit
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/array_obj_ref_232_Merge/merge_req
      -- CP-element group 167: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_232_Update/$exit
      -- 
    ca_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_232_load_0_ack_1, ack => dotP_odd_CP_995_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	18 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/word_0/rr
      -- CP-element group 168: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/word_0/$entry
      -- CP-element group 168: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/$entry
      -- 
    rr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(168), ack => array_obj_ref_236_load_0_req_0); -- 
    dotP_odd_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(170);
      gj_dotP_odd_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	12 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/$entry
      -- CP-element group 169: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/word_0/cr
      -- CP-element group 169: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/word_0/$entry
      -- CP-element group 169: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_update_start_
      -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(169), ack => array_obj_ref_236_load_0_req_1); -- 
    dotP_odd_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(171);
      gj_dotP_odd_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: 	16 
    -- CP-element group 170:  members (5) 
      -- CP-element group 170: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/word_0/ra
      -- CP-element group 170: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/word_0/$exit
      -- CP-element group 170: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Sample/word_access_start/$exit
      -- CP-element group 170: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_sample_completed_
      -- 
    ra_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_236_load_0_ack_0, ack => dotP_odd_CP_995_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	197 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	70 
    -- CP-element group 171:  members (9) 
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/word_0/$exit
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/$exit
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/array_obj_ref_236_Merge/$entry
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/word_access_complete/word_0/ca
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/array_obj_ref_236_Merge/merge_req
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/array_obj_ref_236_Merge/merge_ack
      -- CP-element group 171: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_236_Update/array_obj_ref_236_Merge/$exit
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_236_load_0_ack_1, ack => dotP_odd_CP_995_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	18 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (5) 
      -- CP-element group 172: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/$entry
      -- CP-element group 172: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/word_0/rr
      -- CP-element group 172: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/word_0/$entry
      -- 
    rr_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(172), ack => array_obj_ref_240_load_0_req_0); -- 
    dotP_odd_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(174);
      gj_dotP_odd_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	12 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_update_start_
      -- CP-element group 173: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/word_0/cr
      -- CP-element group 173: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/word_0/$entry
      -- CP-element group 173: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/$entry
      -- 
    cr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(173), ack => array_obj_ref_240_load_0_req_1); -- 
    dotP_odd_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(175);
      gj_dotP_odd_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	16 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/word_0/ra
      -- CP-element group 174: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/$exit
      -- CP-element group 174: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Sample/word_access_start/word_0/$exit
      -- 
    ra_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_240_load_0_ack_0, ack => dotP_odd_CP_995_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	197 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	89 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/array_obj_ref_240_Merge/merge_ack
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/array_obj_ref_240_Merge/merge_req
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/array_obj_ref_240_Merge/$exit
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/array_obj_ref_240_Merge/$entry
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/word_0/ca
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/word_0/$exit
      -- CP-element group 175: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/array_obj_ref_240_Update/word_access_complete/$exit
      -- 
    ca_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_240_load_0_ack_1, ack => dotP_odd_CP_995_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	37 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Sample/req
      -- CP-element group 176: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_sample_start_
      -- 
    req_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(176), ack => W_val_0_231_delayed_5_0_242_inst_req_0); -- 
    dotP_odd_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(37) & dotP_odd_CP_995_elements(178);
      gj_dotP_odd_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	12 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Update/req
      -- CP-element group 177: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_update_start_
      -- 
    req_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(177), ack => W_val_0_231_delayed_5_0_242_inst_req_1); -- 
    dotP_odd_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(179);
      gj_dotP_odd_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	33 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Sample/ack
      -- CP-element group 178: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_sample_completed_
      -- 
    ack_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_0_231_delayed_5_0_242_inst_ack_0, ack => dotP_odd_CP_995_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	197 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	32 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Update/ack
      -- CP-element group 179: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_244_update_completed_
      -- 
    ack_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_0_231_delayed_5_0_242_inst_ack_1, ack => dotP_odd_CP_995_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	56 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Sample/req
      -- CP-element group 180: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_sample_start_
      -- 
    req_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(180), ack => W_val_1_243_delayed_5_0_257_inst_req_0); -- 
    dotP_odd_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(56) & dotP_odd_CP_995_elements(182);
      gj_dotP_odd_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	12 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Update/req
      -- CP-element group 181: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_update_start_
      -- 
    req_1919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(181), ack => W_val_1_243_delayed_5_0_257_inst_req_1); -- 
    dotP_odd_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(183);
      gj_dotP_odd_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: 	52 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Sample/ack
      -- CP-element group 182: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_sample_completed_
      -- 
    ack_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_1_243_delayed_5_0_257_inst_ack_0, ack => dotP_odd_CP_995_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	197 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: 	51 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Update/ack
      -- CP-element group 183: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_259_update_completed_
      -- 
    ack_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_1_243_delayed_5_0_257_inst_ack_1, ack => dotP_odd_CP_995_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	75 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Sample/req
      -- CP-element group 184: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Sample/$entry
      -- 
    req_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(184), ack => W_val_2_255_delayed_5_0_272_inst_req_0); -- 
    dotP_odd_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(75) & dotP_odd_CP_995_elements(186);
      gj_dotP_odd_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	12 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Update/req
      -- CP-element group 185: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_update_start_
      -- 
    req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(185), ack => W_val_2_255_delayed_5_0_272_inst_req_1); -- 
    dotP_odd_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(187);
      gj_dotP_odd_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	71 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Sample/ack
      -- 
    ack_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_2_255_delayed_5_0_272_inst_ack_0, ack => dotP_odd_CP_995_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	197 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	70 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Update/ack
      -- CP-element group 187: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_274_update_completed_
      -- 
    ack_1934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_2_255_delayed_5_0_272_inst_ack_1, ack => dotP_odd_CP_995_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	94 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Sample/req
      -- 
    req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(188), ack => W_val_3_267_delayed_5_0_287_inst_req_0); -- 
    dotP_odd_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(94) & dotP_odd_CP_995_elements(190);
      gj_dotP_odd_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	12 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Update/req
      -- CP-element group 189: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_update_start_
      -- CP-element group 189: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Update/$entry
      -- 
    req_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(189), ack => W_val_3_267_delayed_5_0_287_inst_req_1); -- 
    dotP_odd_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(191);
      gj_dotP_odd_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: 	90 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Sample/ack
      -- CP-element group 190: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Sample/$exit
      -- 
    ack_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_3_267_delayed_5_0_287_inst_ack_0, ack => dotP_odd_CP_995_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	197 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	89 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Update/ack
      -- CP-element group 191: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/assign_stmt_289_update_completed_
      -- 
    ack_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_val_3_267_delayed_5_0_287_inst_ack_1, ack => dotP_odd_CP_995_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	18 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Sample/$entry
      -- 
    rr_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(192), ack => ADD_u8_u8_305_inst_req_0); -- 
    dotP_odd_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(18) & dotP_odd_CP_995_elements(194);
      gj_dotP_odd_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	12 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_update_start_
      -- CP-element group 193: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Update/cr
      -- CP-element group 193: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Update/$entry
      -- 
    cr_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => dotP_odd_CP_995_elements(193), ack => ADD_u8_u8_305_inst_req_1); -- 
    dotP_odd_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(12) & dotP_odd_CP_995_elements(195);
      gj_dotP_odd_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	16 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Sample/ra
      -- 
    ra_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_305_inst_ack_0, ack => dotP_odd_CP_995_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	10 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	15 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/ADD_u8_u8_305_Update/ca
      -- 
    ca_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_305_inst_ack_1, ack => dotP_odd_CP_995_elements(195)); -- 
    -- CP-element group 196:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	9 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	10 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group dotP_odd_CP_995_elements(196) is a control-delay.
    cp_element_196_delay: control_delay_element  generic map(name => " 196_delay", delay_value => 1)  port map(req => dotP_odd_CP_995_elements(9), ack => dotP_odd_CP_995_elements(196), clk => clk, reset =>reset);
    -- CP-element group 197:  join  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	171 
    -- CP-element group 197: 	163 
    -- CP-element group 197: 	167 
    -- CP-element group 197: 	179 
    -- CP-element group 197: 	183 
    -- CP-element group 197: 	156 
    -- CP-element group 197: 	146 
    -- CP-element group 197: 	143 
    -- CP-element group 197: 	139 
    -- CP-element group 197: 	126 
    -- CP-element group 197: 	133 
    -- CP-element group 197: 	130 
    -- CP-element group 197: 	175 
    -- CP-element group 197: 	152 
    -- CP-element group 197: 	187 
    -- CP-element group 197: 	191 
    -- CP-element group 197: 	159 
    -- CP-element group 197: 	113 
    -- CP-element group 197: 	117 
    -- CP-element group 197: 	120 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	6 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_173/do_while_stmt_174/do_while_stmt_174_loop_body/$exit
      -- 
    dotP_odd_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 19) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15);
      constant place_markings: IntegerArray(0 to 19)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant place_delays: IntegerArray(0 to 19) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant joinName: string(1 to 29) := "dotP_odd_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 20); -- 
    begin -- 
      preds <= dotP_odd_CP_995_elements(171) & dotP_odd_CP_995_elements(163) & dotP_odd_CP_995_elements(167) & dotP_odd_CP_995_elements(179) & dotP_odd_CP_995_elements(183) & dotP_odd_CP_995_elements(156) & dotP_odd_CP_995_elements(146) & dotP_odd_CP_995_elements(143) & dotP_odd_CP_995_elements(139) & dotP_odd_CP_995_elements(126) & dotP_odd_CP_995_elements(133) & dotP_odd_CP_995_elements(130) & dotP_odd_CP_995_elements(175) & dotP_odd_CP_995_elements(152) & dotP_odd_CP_995_elements(187) & dotP_odd_CP_995_elements(191) & dotP_odd_CP_995_elements(159) & dotP_odd_CP_995_elements(113) & dotP_odd_CP_995_elements(117) & dotP_odd_CP_995_elements(120);
      gj_dotP_odd_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 20, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => dotP_odd_CP_995_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	5 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_173/do_while_stmt_174/loop_exit/ack
      -- CP-element group 198: 	 branch_block_stmt_173/do_while_stmt_174/loop_exit/$exit
      -- 
    ack_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_174_branch_ack_0, ack => dotP_odd_CP_995_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	5 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_173/do_while_stmt_174/loop_taken/$exit
      -- CP-element group 199: 	 branch_block_stmt_173/do_while_stmt_174/loop_taken/ack
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_174_branch_ack_1, ack => dotP_odd_CP_995_elements(199)); -- 
    -- CP-element group 200:  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	3 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	1 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_173/do_while_stmt_174/$exit
      -- 
    dotP_odd_CP_995_elements(200) <= dotP_odd_CP_995_elements(3);
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	1 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_320/ADD_u32_u32_319_sample_completed_
      -- CP-element group 201: 	 assign_stmt_320/ADD_u32_u32_319_Sample/ra
      -- CP-element group 201: 	 assign_stmt_320/ADD_u32_u32_319_Sample/$exit
      -- 
    ra_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_319_inst_ack_0, ack => dotP_odd_CP_995_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	1 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (5) 
      -- CP-element group 202: 	 assign_stmt_320/ADD_u32_u32_319_update_completed_
      -- CP-element group 202: 	 assign_stmt_320/$exit
      -- CP-element group 202: 	 $exit
      -- CP-element group 202: 	 assign_stmt_320/ADD_u32_u32_319_Update/ca
      -- CP-element group 202: 	 assign_stmt_320/ADD_u32_u32_319_Update/$exit
      -- 
    ca_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_319_inst_ack_1, ack => dotP_odd_CP_995_elements(202)); -- 
    dotP_odd_do_while_stmt_174_terminator_1972: loop_terminator -- 
      generic map (name => " dotP_odd_do_while_stmt_174_terminator_1972", max_iterations_in_flight =>15) 
      port map(loop_body_exit => dotP_odd_CP_995_elements(6),loop_continue => dotP_odd_CP_995_elements(199),loop_terminate => dotP_odd_CP_995_elements(198),loop_back => dotP_odd_CP_995_elements(4),loop_exit => dotP_odd_CP_995_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_176_phi_seq_1068_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_odd_CP_995_elements(21);
      dotP_odd_CP_995_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_odd_CP_995_elements(24);
      dotP_odd_CP_995_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_odd_CP_995_elements(26);
      dotP_odd_CP_995_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_odd_CP_995_elements(19);
      dotP_odd_CP_995_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_odd_CP_995_elements(30);
      dotP_odd_CP_995_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_odd_CP_995_elements(31);
      dotP_odd_CP_995_elements(20) <= phi_mux_reqs(1);
      phi_stmt_176_phi_seq_1068 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_176_phi_seq_1068") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_odd_CP_995_elements(11), 
          phi_sample_ack => dotP_odd_CP_995_elements(17), 
          phi_update_req => dotP_odd_CP_995_elements(13), 
          phi_update_ack => dotP_odd_CP_995_elements(18), 
          phi_mux_ack => dotP_odd_CP_995_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_181_phi_seq_1112_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_odd_CP_995_elements(40);
      dotP_odd_CP_995_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_odd_CP_995_elements(43);
      dotP_odd_CP_995_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_odd_CP_995_elements(45);
      dotP_odd_CP_995_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_odd_CP_995_elements(38);
      dotP_odd_CP_995_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_odd_CP_995_elements(49);
      dotP_odd_CP_995_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_odd_CP_995_elements(50);
      dotP_odd_CP_995_elements(39) <= phi_mux_reqs(1);
      phi_stmt_181_phi_seq_1112 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_181_phi_seq_1112") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_odd_CP_995_elements(34), 
          phi_sample_ack => dotP_odd_CP_995_elements(35), 
          phi_update_req => dotP_odd_CP_995_elements(36), 
          phi_update_ack => dotP_odd_CP_995_elements(37), 
          phi_mux_ack => dotP_odd_CP_995_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_186_phi_seq_1156_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_odd_CP_995_elements(59);
      dotP_odd_CP_995_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_odd_CP_995_elements(62);
      dotP_odd_CP_995_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_odd_CP_995_elements(64);
      dotP_odd_CP_995_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_odd_CP_995_elements(57);
      dotP_odd_CP_995_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_odd_CP_995_elements(68);
      dotP_odd_CP_995_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_odd_CP_995_elements(69);
      dotP_odd_CP_995_elements(58) <= phi_mux_reqs(1);
      phi_stmt_186_phi_seq_1156 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_186_phi_seq_1156") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_odd_CP_995_elements(53), 
          phi_sample_ack => dotP_odd_CP_995_elements(54), 
          phi_update_req => dotP_odd_CP_995_elements(55), 
          phi_update_ack => dotP_odd_CP_995_elements(56), 
          phi_mux_ack => dotP_odd_CP_995_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_191_phi_seq_1200_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_odd_CP_995_elements(78);
      dotP_odd_CP_995_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_odd_CP_995_elements(81);
      dotP_odd_CP_995_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_odd_CP_995_elements(83);
      dotP_odd_CP_995_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_odd_CP_995_elements(76);
      dotP_odd_CP_995_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_odd_CP_995_elements(87);
      dotP_odd_CP_995_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_odd_CP_995_elements(88);
      dotP_odd_CP_995_elements(77) <= phi_mux_reqs(1);
      phi_stmt_191_phi_seq_1200 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_191_phi_seq_1200") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_odd_CP_995_elements(72), 
          phi_sample_ack => dotP_odd_CP_995_elements(73), 
          phi_update_req => dotP_odd_CP_995_elements(74), 
          phi_update_ack => dotP_odd_CP_995_elements(75), 
          phi_mux_ack => dotP_odd_CP_995_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_196_phi_seq_1244_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= dotP_odd_CP_995_elements(97);
      dotP_odd_CP_995_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= dotP_odd_CP_995_elements(100);
      dotP_odd_CP_995_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= dotP_odd_CP_995_elements(102);
      dotP_odd_CP_995_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= dotP_odd_CP_995_elements(95);
      dotP_odd_CP_995_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= dotP_odd_CP_995_elements(106);
      dotP_odd_CP_995_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= dotP_odd_CP_995_elements(107);
      dotP_odd_CP_995_elements(96) <= phi_mux_reqs(1);
      phi_stmt_196_phi_seq_1244 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_196_phi_seq_1244") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => dotP_odd_CP_995_elements(91), 
          phi_sample_ack => dotP_odd_CP_995_elements(92), 
          phi_update_req => dotP_odd_CP_995_elements(93), 
          phi_update_ack => dotP_odd_CP_995_elements(94), 
          phi_mux_ack => dotP_odd_CP_995_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1020_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= dotP_odd_CP_995_elements(7);
        preds(1)  <= dotP_odd_CP_995_elements(8);
        entry_tmerge_1020 : transition_merge -- 
          generic map(name => " entry_tmerge_1020")
          port map (preds => preds, symbol_out => dotP_odd_CP_995_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_317_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_318_wire : std_logic_vector(31 downto 0);
    signal C_176 : std_logic_vector(7 downto 0);
    signal Cr_205 : std_logic_vector(5 downto 0);
    signal MUL_u32_u32_249_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_264_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_279_wire : std_logic_vector(31 downto 0);
    signal MUL_u32_u32_294_wire : std_logic_vector(31 downto 0);
    signal R_Cr_208_resized : std_logic_vector(7 downto 0);
    signal R_Cr_208_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_213_resized : std_logic_vector(7 downto 0);
    signal R_Cr_213_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_218_resized : std_logic_vector(7 downto 0);
    signal R_Cr_218_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_223_resized : std_logic_vector(7 downto 0);
    signal R_Cr_223_scaled : std_logic_vector(7 downto 0);
    signal R_Cr_227_resized : std_logic_vector(2 downto 0);
    signal R_Cr_227_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_231_resized : std_logic_vector(2 downto 0);
    signal R_Cr_231_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_235_resized : std_logic_vector(2 downto 0);
    signal R_Cr_235_scaled : std_logic_vector(2 downto 0);
    signal R_Cr_239_resized : std_logic_vector(2 downto 0);
    signal R_Cr_239_scaled : std_logic_vector(2 downto 0);
    signal R_R_207_resized : std_logic_vector(7 downto 0);
    signal R_R_207_scaled : std_logic_vector(7 downto 0);
    signal R_R_212_resized : std_logic_vector(7 downto 0);
    signal R_R_212_scaled : std_logic_vector(7 downto 0);
    signal R_R_217_resized : std_logic_vector(7 downto 0);
    signal R_R_217_scaled : std_logic_vector(7 downto 0);
    signal R_R_222_resized : std_logic_vector(7 downto 0);
    signal R_R_222_scaled : std_logic_vector(7 downto 0);
    signal ULT_u8_u1_310_wire : std_logic_vector(0 downto 0);
    signal a_rc_0_210 : std_logic_vector(31 downto 0);
    signal a_rc_1_215 : std_logic_vector(31 downto 0);
    signal a_rc_2_220 : std_logic_vector(31 downto 0);
    signal a_rc_3_225 : std_logic_vector(31 downto 0);
    signal array_obj_ref_209_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_209_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_209_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_214_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_214_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_219_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_219_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_224_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_224_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_228_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_228_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_228_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_228_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_228_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_228_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_228_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_232_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_232_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_236_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_236_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_240_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_240_word_offset_0 : std_logic_vector(2 downto 0);
    signal konst_304_wire_constant : std_logic_vector(7 downto 0);
    signal konst_309_wire_constant : std_logic_vector(7 downto 0);
    signal nC_306 : std_logic_vector(7 downto 0);
    signal nC_306_180_buffered : std_logic_vector(7 downto 0);
    signal nval_0_251 : std_logic_vector(31 downto 0);
    signal nval_0_251_185_buffered : std_logic_vector(31 downto 0);
    signal nval_1_266 : std_logic_vector(31 downto 0);
    signal nval_1_266_190_buffered : std_logic_vector(31 downto 0);
    signal nval_2_281 : std_logic_vector(31 downto 0);
    signal nval_2_281_195_buffered : std_logic_vector(31 downto 0);
    signal nval_3_296 : std_logic_vector(31 downto 0);
    signal nval_3_296_200_buffered : std_logic_vector(31 downto 0);
    signal type_cast_179_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_184_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_189_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(31 downto 0);
    signal val_0_181 : std_logic_vector(31 downto 0);
    signal val_0_231_delayed_5_0_244 : std_logic_vector(31 downto 0);
    signal val_1_186 : std_logic_vector(31 downto 0);
    signal val_1_243_delayed_5_0_259 : std_logic_vector(31 downto 0);
    signal val_2_191 : std_logic_vector(31 downto 0);
    signal val_2_255_delayed_5_0_274 : std_logic_vector(31 downto 0);
    signal val_3_196 : std_logic_vector(31 downto 0);
    signal val_3_267_delayed_5_0_289 : std_logic_vector(31 downto 0);
    signal xval_0_229 : std_logic_vector(31 downto 0);
    signal xval_1_233 : std_logic_vector(31 downto 0);
    signal xval_2_237 : std_logic_vector(31 downto 0);
    signal xval_3_241 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_209_offset_scale_factor_0 <= "00001000";
    array_obj_ref_209_offset_scale_factor_1 <= "00000001";
    array_obj_ref_209_resized_base_address <= "00000000";
    array_obj_ref_209_word_offset_0 <= "00000000";
    array_obj_ref_214_offset_scale_factor_0 <= "00001000";
    array_obj_ref_214_offset_scale_factor_1 <= "00000001";
    array_obj_ref_214_resized_base_address <= "00000000";
    array_obj_ref_214_word_offset_0 <= "00000000";
    array_obj_ref_219_offset_scale_factor_0 <= "00001000";
    array_obj_ref_219_offset_scale_factor_1 <= "00000001";
    array_obj_ref_219_resized_base_address <= "00000000";
    array_obj_ref_219_word_offset_0 <= "00000000";
    array_obj_ref_224_offset_scale_factor_0 <= "00001000";
    array_obj_ref_224_offset_scale_factor_1 <= "00000001";
    array_obj_ref_224_resized_base_address <= "00000000";
    array_obj_ref_224_word_offset_0 <= "00000000";
    array_obj_ref_228_offset_scale_factor_0 <= "001";
    array_obj_ref_228_resized_base_address <= "000";
    array_obj_ref_228_word_offset_0 <= "000";
    array_obj_ref_232_offset_scale_factor_0 <= "001";
    array_obj_ref_232_resized_base_address <= "000";
    array_obj_ref_232_word_offset_0 <= "000";
    array_obj_ref_236_offset_scale_factor_0 <= "001";
    array_obj_ref_236_resized_base_address <= "000";
    array_obj_ref_236_word_offset_0 <= "000";
    array_obj_ref_240_offset_scale_factor_0 <= "001";
    array_obj_ref_240_resized_base_address <= "000";
    array_obj_ref_240_word_offset_0 <= "000";
    konst_304_wire_constant <= "00000100";
    konst_309_wire_constant <= "00100000";
    type_cast_179_wire_constant <= "00000000";
    type_cast_184_wire_constant <= "00000000000000000000000000000000";
    type_cast_189_wire_constant <= "00000000000000000000000000000000";
    type_cast_194_wire_constant <= "00000000000000000000000000000000";
    type_cast_199_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_176: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_179_wire_constant & nC_306_180_buffered;
      req <= phi_stmt_176_req_0 & phi_stmt_176_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_176",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_176_ack_0,
          idata => idata,
          odata => C_176,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_176
    phi_stmt_181: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_184_wire_constant & nval_0_251_185_buffered;
      req <= phi_stmt_181_req_0 & phi_stmt_181_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_181",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_181_ack_0,
          idata => idata,
          odata => val_0_181,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_181
    phi_stmt_186: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_189_wire_constant & nval_1_266_190_buffered;
      req <= phi_stmt_186_req_0 & phi_stmt_186_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_186",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_186_ack_0,
          idata => idata,
          odata => val_1_186,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_186
    phi_stmt_191: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_194_wire_constant & nval_2_281_195_buffered;
      req <= phi_stmt_191_req_0 & phi_stmt_191_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_191",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_191_ack_0,
          idata => idata,
          odata => val_2_191,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_191
    phi_stmt_196: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_199_wire_constant & nval_3_296_200_buffered;
      req <= phi_stmt_196_req_0 & phi_stmt_196_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_196",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_196_ack_0,
          idata => idata,
          odata => val_3_196,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_196
    -- flow-through slice operator slice_204_inst
    Cr_205 <= C_176(7 downto 2);
    W_val_0_231_delayed_5_0_242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_0_231_delayed_5_0_242_inst_req_0;
      W_val_0_231_delayed_5_0_242_inst_ack_0<= wack(0);
      rreq(0) <= W_val_0_231_delayed_5_0_242_inst_req_1;
      W_val_0_231_delayed_5_0_242_inst_ack_1<= rack(0);
      W_val_0_231_delayed_5_0_242_inst : InterlockBuffer generic map ( -- 
        name => "W_val_0_231_delayed_5_0_242_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_0_181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_0_231_delayed_5_0_244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_1_243_delayed_5_0_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_1_243_delayed_5_0_257_inst_req_0;
      W_val_1_243_delayed_5_0_257_inst_ack_0<= wack(0);
      rreq(0) <= W_val_1_243_delayed_5_0_257_inst_req_1;
      W_val_1_243_delayed_5_0_257_inst_ack_1<= rack(0);
      W_val_1_243_delayed_5_0_257_inst : InterlockBuffer generic map ( -- 
        name => "W_val_1_243_delayed_5_0_257_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_1_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_1_243_delayed_5_0_259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_2_255_delayed_5_0_272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_2_255_delayed_5_0_272_inst_req_0;
      W_val_2_255_delayed_5_0_272_inst_ack_0<= wack(0);
      rreq(0) <= W_val_2_255_delayed_5_0_272_inst_req_1;
      W_val_2_255_delayed_5_0_272_inst_ack_1<= rack(0);
      W_val_2_255_delayed_5_0_272_inst : InterlockBuffer generic map ( -- 
        name => "W_val_2_255_delayed_5_0_272_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_2_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_2_255_delayed_5_0_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_val_3_267_delayed_5_0_287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_val_3_267_delayed_5_0_287_inst_req_0;
      W_val_3_267_delayed_5_0_287_inst_ack_0<= wack(0);
      rreq(0) <= W_val_3_267_delayed_5_0_287_inst_req_1;
      W_val_3_267_delayed_5_0_287_inst_ack_1<= rack(0);
      W_val_3_267_delayed_5_0_287_inst : InterlockBuffer generic map ( -- 
        name => "W_val_3_267_delayed_5_0_287_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => val_3_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => val_3_267_delayed_5_0_289,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nC_306_180_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nC_306_180_buf_req_0;
      nC_306_180_buf_ack_0<= wack(0);
      rreq(0) <= nC_306_180_buf_req_1;
      nC_306_180_buf_ack_1<= rack(0);
      nC_306_180_buf : InterlockBuffer generic map ( -- 
        name => "nC_306_180_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nC_306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nC_306_180_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_0_251_185_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_0_251_185_buf_req_0;
      nval_0_251_185_buf_ack_0<= wack(0);
      rreq(0) <= nval_0_251_185_buf_req_1;
      nval_0_251_185_buf_ack_1<= rack(0);
      nval_0_251_185_buf : InterlockBuffer generic map ( -- 
        name => "nval_0_251_185_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_0_251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_0_251_185_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_1_266_190_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_1_266_190_buf_req_0;
      nval_1_266_190_buf_ack_0<= wack(0);
      rreq(0) <= nval_1_266_190_buf_req_1;
      nval_1_266_190_buf_ack_1<= rack(0);
      nval_1_266_190_buf : InterlockBuffer generic map ( -- 
        name => "nval_1_266_190_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_1_266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_1_266_190_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_2_281_195_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_2_281_195_buf_req_0;
      nval_2_281_195_buf_ack_0<= wack(0);
      rreq(0) <= nval_2_281_195_buf_req_1;
      nval_2_281_195_buf_ack_1<= rack(0);
      nval_2_281_195_buf : InterlockBuffer generic map ( -- 
        name => "nval_2_281_195_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_2_281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_2_281_195_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nval_3_296_200_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nval_3_296_200_buf_req_0;
      nval_3_296_200_buf_ack_0<= wack(0);
      rreq(0) <= nval_3_296_200_buf_req_1;
      nval_3_296_200_buf_ack_1<= rack(0);
      nval_3_296_200_buf : InterlockBuffer generic map ( -- 
        name => "nval_3_296_200_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nval_3_296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nval_3_296_200_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_209_addr_0
    process(array_obj_ref_209_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_209_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_209_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_gather_scatter
    process(array_obj_ref_209_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_209_data_0;
      ov(31 downto 0) := iv;
      a_rc_0_210 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_207_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_index_1_rename
    process(R_Cr_208_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_208_resized;
      ov(7 downto 0) := iv;
      R_Cr_208_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_index_1_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov(5 downto 0) := iv;
      R_Cr_208_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_index_offset
    process(array_obj_ref_209_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_209_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_209_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_209_root_address_inst
    process(array_obj_ref_209_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_209_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_209_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_addr_0
    process(array_obj_ref_214_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_214_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_214_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_gather_scatter
    process(array_obj_ref_214_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_214_data_0;
      ov(31 downto 0) := iv;
      a_rc_1_215 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_212_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_index_1_rename
    process(R_Cr_213_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_213_resized;
      ov(7 downto 0) := iv;
      R_Cr_213_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_index_1_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov(5 downto 0) := iv;
      R_Cr_213_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_index_offset
    process(array_obj_ref_214_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_214_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_214_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_214_root_address_inst
    process(array_obj_ref_214_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_214_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_214_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_addr_0
    process(array_obj_ref_219_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_219_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_219_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_gather_scatter
    process(array_obj_ref_219_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_219_data_0;
      ov(31 downto 0) := iv;
      a_rc_2_220 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_217_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_index_1_rename
    process(R_Cr_218_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_218_resized;
      ov(7 downto 0) := iv;
      R_Cr_218_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_index_1_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov(5 downto 0) := iv;
      R_Cr_218_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_index_offset
    process(array_obj_ref_219_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_219_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_219_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_219_root_address_inst
    process(array_obj_ref_219_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_219_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_219_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_addr_0
    process(array_obj_ref_224_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_224_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_224_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_gather_scatter
    process(array_obj_ref_224_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_224_data_0;
      ov(31 downto 0) := iv;
      a_rc_3_225 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_index_0_resize
    process(R_buffer) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_buffer;
      ov(7 downto 0) := iv;
      R_R_222_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_index_1_rename
    process(R_Cr_223_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_223_resized;
      ov(7 downto 0) := iv;
      R_Cr_223_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_index_1_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov(5 downto 0) := iv;
      R_Cr_223_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_index_offset
    process(array_obj_ref_224_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_224_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_224_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_224_root_address_inst
    process(array_obj_ref_224_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_224_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_224_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_addr_0
    process(array_obj_ref_228_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_228_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_228_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_gather_scatter
    process(array_obj_ref_228_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_228_data_0;
      ov(31 downto 0) := iv;
      xval_0_229 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_0_rename
    process(R_Cr_227_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_227_resized;
      ov(2 downto 0) := iv;
      R_Cr_227_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_0_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov := iv(2 downto 0);
      R_Cr_227_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_index_offset
    process(R_Cr_227_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_227_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_228_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_228_root_address_inst
    process(array_obj_ref_228_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_228_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_228_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_addr_0
    process(array_obj_ref_232_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_232_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_232_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_gather_scatter
    process(array_obj_ref_232_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_232_data_0;
      ov(31 downto 0) := iv;
      xval_1_233 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_index_0_rename
    process(R_Cr_231_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_231_resized;
      ov(2 downto 0) := iv;
      R_Cr_231_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_index_0_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov := iv(2 downto 0);
      R_Cr_231_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_index_offset
    process(R_Cr_231_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_231_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_232_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_232_root_address_inst
    process(array_obj_ref_232_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_232_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_232_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_addr_0
    process(array_obj_ref_236_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_236_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_236_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_gather_scatter
    process(array_obj_ref_236_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_236_data_0;
      ov(31 downto 0) := iv;
      xval_2_237 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_index_0_rename
    process(R_Cr_235_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_235_resized;
      ov(2 downto 0) := iv;
      R_Cr_235_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_index_0_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov := iv(2 downto 0);
      R_Cr_235_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_index_offset
    process(R_Cr_235_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_235_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_236_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_236_root_address_inst
    process(array_obj_ref_236_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_236_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_236_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_addr_0
    process(array_obj_ref_240_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_240_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_240_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_gather_scatter
    process(array_obj_ref_240_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_240_data_0;
      ov(31 downto 0) := iv;
      xval_3_241 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_index_0_rename
    process(R_Cr_239_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_239_resized;
      ov(2 downto 0) := iv;
      R_Cr_239_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_index_0_resize
    process(Cr_205) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Cr_205;
      ov := iv(2 downto 0);
      R_Cr_239_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_index_offset
    process(R_Cr_239_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Cr_239_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_240_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_240_root_address_inst
    process(array_obj_ref_240_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_240_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_240_root_address <= ov(2 downto 0);
      --
    end process;
    do_while_stmt_174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_310_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_174_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_174_branch_req_0,
          ack0 => do_while_stmt_174_branch_ack_0,
          ack1 => do_while_stmt_174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_250_inst
    process(val_0_231_delayed_5_0_244, MUL_u32_u32_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_0_231_delayed_5_0_244, MUL_u32_u32_249_wire, tmp_var);
      nval_0_251 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_265_inst
    process(val_1_243_delayed_5_0_259, MUL_u32_u32_264_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_1_243_delayed_5_0_259, MUL_u32_u32_264_wire, tmp_var);
      nval_1_266 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_280_inst
    process(val_2_255_delayed_5_0_274, MUL_u32_u32_279_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_2_255_delayed_5_0_274, MUL_u32_u32_279_wire, tmp_var);
      nval_2_281 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_295_inst
    process(val_3_267_delayed_5_0_289, MUL_u32_u32_294_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(val_3_267_delayed_5_0_289, MUL_u32_u32_294_wire, tmp_var);
      nval_3_296 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_317_inst
    process(nval_2_281, nval_3_296) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nval_2_281, nval_3_296, tmp_var);
      ADD_u32_u32_317_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_318_inst
    process(nval_1_266, ADD_u32_u32_317_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nval_1_266, ADD_u32_u32_317_wire, tmp_var);
      ADD_u32_u32_318_wire <= tmp_var; --
    end process;
    -- shared split operator group (6) : ADD_u32_u32_319_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= nval_0_251 & ADD_u32_u32_318_wire;
      result_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_319_inst_req_0;
      ADD_u32_u32_319_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_319_inst_req_1;
      ADD_u32_u32_319_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : ADD_u8_u8_305_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= C_176;
      nC_306 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_305_inst_req_0;
      ADD_u8_u8_305_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_305_inst_req_1;
      ADD_u8_u8_305_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000100",
          constant_width => 8,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator MUL_u32_u32_249_inst
    process(a_rc_0_210, xval_0_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_0_210, xval_0_229, tmp_var);
      MUL_u32_u32_249_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_264_inst
    process(a_rc_1_215, xval_1_233) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_1_215, xval_1_233, tmp_var);
      MUL_u32_u32_264_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_279_inst
    process(a_rc_2_220, xval_2_237) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_2_220, xval_2_237, tmp_var);
      MUL_u32_u32_279_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_294_inst
    process(a_rc_3_225, xval_3_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(a_rc_3_225, xval_3_241, tmp_var);
      MUL_u32_u32_294_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_310_inst
    process(nC_306) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nC_306, konst_309_wire_constant, tmp_var);
      ULT_u8_u1_310_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_209_index_0_scale array_obj_ref_214_index_0_scale array_obj_ref_219_index_0_scale array_obj_ref_224_index_0_scale 
    ApIntMul_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      data_in <= R_R_207_resized & R_R_212_resized & R_R_217_resized & R_R_222_resized;
      R_R_207_scaled <= data_out(31 downto 24);
      R_R_212_scaled <= data_out(23 downto 16);
      R_R_217_scaled <= data_out(15 downto 8);
      R_R_222_scaled <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      reqL_unguarded(3) <= array_obj_ref_209_index_0_scale_req_0;
      reqL_unguarded(2) <= array_obj_ref_214_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_219_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_224_index_0_scale_req_0;
      array_obj_ref_209_index_0_scale_ack_0 <= ackL_unguarded(3);
      array_obj_ref_214_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_219_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_224_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_209_index_0_scale_req_1;
      reqR_unguarded(2) <= array_obj_ref_214_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_219_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_224_index_0_scale_req_1;
      array_obj_ref_209_index_0_scale_ack_1 <= ackR_unguarded(3);
      array_obj_ref_214_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_219_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_224_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_13_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_2: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_accessRegulator_3: access_regulator_base generic map (name => "ApIntMul_group_13_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApIntMul_group_13_gI: SplitGuardInterface generic map(name => "ApIntMul_group_13_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_13",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00001000",
          constant_width => 8,
          use_constant  => true,
          full_rate  => true,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 4,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_209_index_sum_1 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_208_scaled & R_R_207_scaled;
      array_obj_ref_209_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_209_index_sum_1_req_0;
      array_obj_ref_209_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_209_index_sum_1_req_1;
      array_obj_ref_209_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_214_index_sum_1 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_213_scaled & R_R_212_scaled;
      array_obj_ref_214_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_214_index_sum_1_req_0;
      array_obj_ref_214_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_214_index_sum_1_req_1;
      array_obj_ref_214_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : array_obj_ref_219_index_sum_1 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_218_scaled & R_R_217_scaled;
      array_obj_ref_219_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_219_index_sum_1_req_0;
      array_obj_ref_219_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_219_index_sum_1_req_1;
      array_obj_ref_219_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : array_obj_ref_224_index_sum_1 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Cr_223_scaled & R_R_222_scaled;
      array_obj_ref_224_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_224_index_sum_1_req_0;
      array_obj_ref_224_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_224_index_sum_1_req_1;
      array_obj_ref_224_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : array_obj_ref_209_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_209_load_0_req_0;
      array_obj_ref_209_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_209_load_0_req_1;
      array_obj_ref_209_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_209_word_address_0;
      array_obj_ref_209_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(7 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : array_obj_ref_214_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_214_load_0_req_0;
      array_obj_ref_214_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_214_load_0_req_1;
      array_obj_ref_214_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_214_word_address_0;
      array_obj_ref_214_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(7 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : array_obj_ref_219_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_219_load_0_req_0;
      array_obj_ref_219_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_219_load_0_req_1;
      array_obj_ref_219_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_219_word_address_0;
      array_obj_ref_219_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(7 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : array_obj_ref_224_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_224_load_0_req_0;
      array_obj_ref_224_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_224_load_0_req_1;
      array_obj_ref_224_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_224_word_address_0;
      array_obj_ref_224_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(7 downto 0),
          mtag => memory_space_3_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : array_obj_ref_228_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_228_load_0_req_0;
      array_obj_ref_228_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_228_load_0_req_1;
      array_obj_ref_228_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_228_word_address_0;
      array_obj_ref_228_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(2 downto 0),
          mtag => memory_space_4_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : array_obj_ref_232_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_232_load_0_req_0;
      array_obj_ref_232_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_232_load_0_req_1;
      array_obj_ref_232_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_232_word_address_0;
      array_obj_ref_232_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(2 downto 0),
          mtag => memory_space_5_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : array_obj_ref_236_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_236_load_0_req_0;
      array_obj_ref_236_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_236_load_0_req_1;
      array_obj_ref_236_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_236_word_address_0;
      array_obj_ref_236_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(2 downto 0),
          mtag => memory_space_6_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : array_obj_ref_240_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_240_load_0_req_0;
      array_obj_ref_240_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_240_load_0_req_1;
      array_obj_ref_240_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup7_gI: SplitGuardInterface generic map(name => "LoadGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_240_word_address_0;
      array_obj_ref_240_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup7", addr_width => 3,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(2 downto 0),
          mtag => memory_space_7_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup7 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(31 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- 
  end Block; -- data_path
  -- 
end dotP_odd_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity multiplyMatrixVector is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
    dotP_even_call_reqs : out  std_logic_vector(0 downto 0);
    dotP_even_call_acks : in   std_logic_vector(0 downto 0);
    dotP_even_call_data : out  std_logic_vector(7 downto 0);
    dotP_even_call_tag  :  out  std_logic_vector(0 downto 0);
    dotP_even_return_reqs : out  std_logic_vector(0 downto 0);
    dotP_even_return_acks : in   std_logic_vector(0 downto 0);
    dotP_even_return_data : in   std_logic_vector(31 downto 0);
    dotP_even_return_tag :  in   std_logic_vector(0 downto 0);
    dotP_odd_call_reqs : out  std_logic_vector(0 downto 0);
    dotP_odd_call_acks : in   std_logic_vector(0 downto 0);
    dotP_odd_call_data : out  std_logic_vector(7 downto 0);
    dotP_odd_call_tag  :  out  std_logic_vector(0 downto 0);
    dotP_odd_return_reqs : out  std_logic_vector(0 downto 0);
    dotP_odd_return_acks : in   std_logic_vector(0 downto 0);
    dotP_odd_return_data : in   std_logic_vector(31 downto 0);
    dotP_odd_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity multiplyMatrixVector;
architecture multiplyMatrixVector_arch of multiplyMatrixVector is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal multiplyMatrixVector_CP_1993_start: Boolean;
  signal multiplyMatrixVector_CP_1993_symbol: Boolean;
  -- volatile/operator module components. 
  component dotP_even is -- 
    generic (tag_length : integer); 
    port ( -- 
      R : in  std_logic_vector(7 downto 0);
      result : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component dotP_odd is -- 
    generic (tag_length : integer); 
    port ( -- 
      R : in  std_logic_vector(7 downto 0);
      result : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_341_call_ack_0 : boolean;
  signal call_stmt_341_call_req_0 : boolean;
  signal call_stmt_336_call_ack_1 : boolean;
  signal call_stmt_336_call_req_1 : boolean;
  signal call_stmt_341_call_ack_1 : boolean;
  signal call_stmt_341_call_req_1 : boolean;
  signal call_stmt_336_call_ack_0 : boolean;
  signal call_stmt_336_call_req_0 : boolean;
  signal array_obj_ref_343_store_0_req_0 : boolean;
  signal array_obj_ref_343_store_0_ack_0 : boolean;
  signal array_obj_ref_343_store_0_req_1 : boolean;
  signal array_obj_ref_343_store_0_ack_1 : boolean;
  signal array_obj_ref_349_store_0_req_0 : boolean;
  signal array_obj_ref_349_store_0_ack_0 : boolean;
  signal array_obj_ref_349_store_0_req_1 : boolean;
  signal array_obj_ref_349_store_0_ack_1 : boolean;
  signal ADD_u8_u8_355_inst_req_0 : boolean;
  signal ADD_u8_u8_355_inst_ack_0 : boolean;
  signal ADD_u8_u8_355_inst_req_1 : boolean;
  signal ADD_u8_u8_355_inst_ack_1 : boolean;
  signal if_stmt_357_branch_req_0 : boolean;
  signal if_stmt_357_branch_ack_1 : boolean;
  signal if_stmt_357_branch_ack_0 : boolean;
  signal phi_stmt_328_req_0 : boolean;
  signal nR_356_332_buf_req_0 : boolean;
  signal nR_356_332_buf_ack_0 : boolean;
  signal nR_356_332_buf_req_1 : boolean;
  signal nR_356_332_buf_ack_1 : boolean;
  signal phi_stmt_328_req_1 : boolean;
  signal phi_stmt_328_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "multiplyMatrixVector_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  multiplyMatrixVector_CP_1993_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "multiplyMatrixVector_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= multiplyMatrixVector_CP_1993_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= multiplyMatrixVector_CP_1993_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= multiplyMatrixVector_CP_1993_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  multiplyMatrixVector_CP_1993: Block -- control-path 
    signal multiplyMatrixVector_CP_1993_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    multiplyMatrixVector_CP_1993_elements(0) <= multiplyMatrixVector_CP_1993_start;
    multiplyMatrixVector_CP_1993_symbol <= multiplyMatrixVector_CP_1993_elements(16);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_326/$entry
      -- CP-element group 0: 	 branch_block_stmt_326/merge_stmt_327__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_326/branch_block_stmt_326__entry__
      -- CP-element group 0: 	 branch_block_stmt_326/merge_stmt_327_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/$entry
      -- CP-element group 0: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/phi_stmt_328_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	22 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Sample/$exit
      -- 
    cra_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_336_call_ack_0, ack => multiplyMatrixVector_CP_1993_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	22 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_update_completed_
      -- 
    cca_2023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_336_call_ack_1, ack => multiplyMatrixVector_CP_1993_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	22 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_sample_completed_
      -- 
    cra_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_341_call_ack_0, ack => multiplyMatrixVector_CP_1993_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	22 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	8 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_update_completed_
      -- 
    cca_2037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_341_call_ack_1, ack => multiplyMatrixVector_CP_1993_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	22 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/array_obj_ref_343_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/array_obj_ref_343_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/array_obj_ref_343_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/array_obj_ref_343_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/word_0/rr
      -- 
    rr_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(5), ack => array_obj_ref_343_store_0_req_0); -- 
    multiplyMatrixVector_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "multiplyMatrixVector_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= multiplyMatrixVector_CP_1993_elements(2) & multiplyMatrixVector_CP_1993_elements(22);
      gj_multiplyMatrixVector_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => multiplyMatrixVector_CP_1993_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	13 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Sample/word_access_start/word_0/ra
      -- 
    ra_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_343_store_0_ack_0, ack => multiplyMatrixVector_CP_1993_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	22 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	14 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/word_0/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_343_store_0_ack_1, ack => multiplyMatrixVector_CP_1993_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	13 
    -- CP-element group 8: 	22 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/array_obj_ref_349_Split/$entry
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/array_obj_ref_349_Split/$exit
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/array_obj_ref_349_Split/split_req
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/array_obj_ref_349_Split/split_ack
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/word_0/rr
      -- 
    rr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(8), ack => array_obj_ref_349_store_0_req_0); -- 
    multiplyMatrixVector_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "multiplyMatrixVector_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= multiplyMatrixVector_CP_1993_elements(4) & multiplyMatrixVector_CP_1993_elements(13) & multiplyMatrixVector_CP_1993_elements(22);
      gj_multiplyMatrixVector_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => multiplyMatrixVector_CP_1993_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Sample/word_access_start/word_0/ra
      -- 
    ra_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_store_0_ack_0, ack => multiplyMatrixVector_CP_1993_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	22 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	14 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/word_0/ca
      -- 
    ca_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_store_0_ack_1, ack => multiplyMatrixVector_CP_1993_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	22 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Sample/ra
      -- 
    ra_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_355_inst_ack_0, ack => multiplyMatrixVector_CP_1993_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	22 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Update/ca
      -- 
    ca_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_355_inst_ack_1, ack => multiplyMatrixVector_CP_1993_elements(12)); -- 
    -- CP-element group 13:  transition  delay-element  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	6 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_array_obj_ref_349_delay
      -- 
    -- Element group multiplyMatrixVector_CP_1993_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => multiplyMatrixVector_CP_1993_elements(6), ack => multiplyMatrixVector_CP_1993_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  branch  join  transition  place  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	7 
    -- CP-element group 14: 	10 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (24) 
      -- CP-element group 14: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356__exit__
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357__entry__
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_dead_link/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/ULT_u8_u1_360_inputs/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/ULT_u8_u1_360_inputs/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/ULT_u8_u1_360/SplitProtocol/Update/ca
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_eval_test/branch_req
      -- CP-element group 14: 	 branch_block_stmt_326/ULT_u8_u1_360_place
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_if_link/$entry
      -- CP-element group 14: 	 branch_block_stmt_326/if_stmt_357_else_link/$entry
      -- 
    branch_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(14), ack => if_stmt_357_branch_req_0); -- 
    multiplyMatrixVector_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "multiplyMatrixVector_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= multiplyMatrixVector_CP_1993_elements(7) & multiplyMatrixVector_CP_1993_elements(10) & multiplyMatrixVector_CP_1993_elements(12);
      gj_multiplyMatrixVector_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => multiplyMatrixVector_CP_1993_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_326/if_stmt_357_if_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_326/if_stmt_357_if_link/if_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_326/loopback
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Sample/req
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Update/req
      -- 
    if_choice_transition_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_357_branch_ack_1, ack => multiplyMatrixVector_CP_1993_elements(15)); -- 
    req_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(15), ack => nR_356_332_buf_req_0); -- 
    req_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(15), ack => nR_356_332_buf_req_1); -- 
    -- CP-element group 16:  merge  transition  place  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_326/$exit
      -- CP-element group 16: 	 branch_block_stmt_326/branch_block_stmt_326__exit__
      -- CP-element group 16: 	 $exit
      -- CP-element group 16: 	 branch_block_stmt_326/if_stmt_357__exit__
      -- CP-element group 16: 	 branch_block_stmt_326/if_stmt_357_else_link/$exit
      -- CP-element group 16: 	 branch_block_stmt_326/if_stmt_357_else_link/else_choice_transition
      -- 
    else_choice_transition_2212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_357_branch_ack_0, ack => multiplyMatrixVector_CP_1993_elements(16)); -- 
    -- CP-element group 17:  transition  output  delay-element  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/$exit
      -- CP-element group 17: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/$exit
      -- CP-element group 17: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/phi_stmt_328_sources/$exit
      -- CP-element group 17: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_331_konst_delay_trans
      -- CP-element group 17: 	 branch_block_stmt_326/merge_stmt_327__entry___PhiReq/phi_stmt_328/phi_stmt_328_req
      -- 
    phi_stmt_328_req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_328_req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(17), ack => phi_stmt_328_req_0); -- 
    -- Element group multiplyMatrixVector_CP_1993_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => multiplyMatrixVector_CP_1993_elements(0), ack => multiplyMatrixVector_CP_1993_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Sample/ack
      -- 
    ack_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_356_332_buf_ack_0, ack => multiplyMatrixVector_CP_1993_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/Update/ack
      -- 
    ack_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_356_332_buf_ack_1, ack => multiplyMatrixVector_CP_1993_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_326/loopback_PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/$exit
      -- CP-element group 20: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/$exit
      -- CP-element group 20: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_sources/Interlock/$exit
      -- CP-element group 20: 	 branch_block_stmt_326/loopback_PhiReq/phi_stmt_328/phi_stmt_328_req
      -- 
    phi_stmt_328_req_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_328_req_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(20), ack => phi_stmt_328_req_1); -- 
    multiplyMatrixVector_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "multiplyMatrixVector_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= multiplyMatrixVector_CP_1993_elements(18) & multiplyMatrixVector_CP_1993_elements(19);
      gj_multiplyMatrixVector_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => multiplyMatrixVector_CP_1993_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  merge  transition  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_326/merge_stmt_327_PhiReqMerge
      -- CP-element group 21: 	 branch_block_stmt_326/merge_stmt_327_PhiAck/$entry
      -- 
    multiplyMatrixVector_CP_1993_elements(21) <= OrReduce(multiplyMatrixVector_CP_1993_elements(17) & multiplyMatrixVector_CP_1993_elements(20));
    -- CP-element group 22:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	1 
    -- CP-element group 22: 	2 
    -- CP-element group 22: 	3 
    -- CP-element group 22: 	4 
    -- CP-element group 22: 	5 
    -- CP-element group 22: 	8 
    -- CP-element group 22: 	7 
    -- CP-element group 22: 	10 
    -- CP-element group 22: 	11 
    -- CP-element group 22: 	12 
    -- CP-element group 22:  members (85) 
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_scale_0/scale_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_326/merge_stmt_327__exit__
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Sample/crr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356__entry__
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_resize_0/index_resize_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_update_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_offset_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Update/ccr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_word_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_root_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Update/ccr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_update_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_resized_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Sample/crr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_336_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_update_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_scale_0/scale_rename_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_base_plus_offset/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_base_plus_offset/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_final_index_sum_regn/ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_computed_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_resize_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_final_index_sum_regn/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_final_index_sum_regn/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_word_addrgen/root_register_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_word_addrgen/root_register_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_scale_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_word_addrgen/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_word_addrgen/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_scaled_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_final_index_sum_regn/req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_resize_0/index_resize_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_scale_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_index_resize_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/call_stmt_341_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/word_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_343_Update/word_access_complete/word_0/cr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_update_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_word_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_root_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_offset_calculated
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_resized_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_scaled_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_computed_0
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_resize_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_resize_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_resize_0/index_resize_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_resize_0/index_resize_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_scale_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_scale_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_scale_0/scale_rename_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_index_scale_0/scale_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_final_index_sum_regn/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_final_index_sum_regn/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_final_index_sum_regn/req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_final_index_sum_regn/ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_base_plus_offset/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_base_plus_offset/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_word_addrgen/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_word_addrgen/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_word_addrgen/root_register_req
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_word_addrgen/root_register_ack
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/word_0/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/array_obj_ref_349_Update/word_access_complete/word_0/cr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_update_start_
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_326/call_stmt_336_to_assign_stmt_356/ADD_u8_u8_355_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_326/merge_stmt_327_PhiAck/$exit
      -- CP-element group 22: 	 branch_block_stmt_326/merge_stmt_327_PhiAck/phi_stmt_328_ack
      -- 
    phi_stmt_328_ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_328_ack_0, ack => multiplyMatrixVector_CP_1993_elements(22)); -- 
    crr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => call_stmt_341_call_req_0); -- 
    ccr_2022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => call_stmt_336_call_req_1); -- 
    ccr_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => call_stmt_341_call_req_1); -- 
    crr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => call_stmt_336_call_req_0); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => array_obj_ref_343_store_0_req_1); -- 
    cr_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => array_obj_ref_349_store_0_req_1); -- 
    rr_2169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => ADD_u8_u8_355_inst_req_0); -- 
    cr_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => multiplyMatrixVector_CP_1993_elements(22), ack => ADD_u8_u8_355_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_339_wire : std_logic_vector(7 downto 0);
    signal ADD_u8_u8_348_resized : std_logic_vector(4 downto 0);
    signal ADD_u8_u8_348_scaled : std_logic_vector(4 downto 0);
    signal ADD_u8_u8_348_wire : std_logic_vector(7 downto 0);
    signal R_328 : std_logic_vector(7 downto 0);
    signal R_R_342_resized : std_logic_vector(4 downto 0);
    signal R_R_342_scaled : std_logic_vector(4 downto 0);
    signal ULT_u8_u1_360_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_343_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_343_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_343_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_343_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_343_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_343_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_343_word_offset_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_349_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_349_word_offset_0 : std_logic_vector(4 downto 0);
    signal konst_338_wire_constant : std_logic_vector(7 downto 0);
    signal konst_347_wire_constant : std_logic_vector(7 downto 0);
    signal konst_354_wire_constant : std_logic_vector(7 downto 0);
    signal konst_359_wire_constant : std_logic_vector(7 downto 0);
    signal nR_356 : std_logic_vector(7 downto 0);
    signal nR_356_332_buffered : std_logic_vector(7 downto 0);
    signal type_cast_331_wire_constant : std_logic_vector(7 downto 0);
    signal val_even_336 : std_logic_vector(31 downto 0);
    signal val_odd_341 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_343_offset_scale_factor_0 <= "00001";
    array_obj_ref_343_resized_base_address <= "00000";
    array_obj_ref_343_word_offset_0 <= "00000";
    array_obj_ref_349_offset_scale_factor_0 <= "00001";
    array_obj_ref_349_resized_base_address <= "00000";
    array_obj_ref_349_word_offset_0 <= "00000";
    konst_338_wire_constant <= "00000001";
    konst_347_wire_constant <= "00000001";
    konst_354_wire_constant <= "00000001";
    konst_359_wire_constant <= "00100000";
    type_cast_331_wire_constant <= "00000000";
    phi_stmt_328: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_331_wire_constant & nR_356_332_buffered;
      req <= phi_stmt_328_req_0 & phi_stmt_328_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_328",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_328_ack_0,
          idata => idata,
          odata => R_328,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_328
    nR_356_332_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_356_332_buf_req_0;
      nR_356_332_buf_ack_0<= wack(0);
      rreq(0) <= nR_356_332_buf_req_1;
      nR_356_332_buf_ack_1<= rack(0);
      nR_356_332_buf : InterlockBuffer generic map ( -- 
        name => "nR_356_332_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_356_332_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_343_addr_0
    process(array_obj_ref_343_root_address) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_343_root_address;
      ov(4 downto 0) := iv;
      array_obj_ref_343_word_address_0 <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_gather_scatter
    process(val_even_336) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_even_336;
      ov(31 downto 0) := iv;
      array_obj_ref_343_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_index_0_rename
    process(R_R_342_resized) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_R_342_resized;
      ov(4 downto 0) := iv;
      R_R_342_scaled <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_index_0_resize
    process(R_328) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_328;
      ov := iv(4 downto 0);
      R_R_342_resized <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_index_offset
    process(R_R_342_scaled) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_R_342_scaled;
      ov(4 downto 0) := iv;
      array_obj_ref_343_final_offset <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_root_address_inst
    process(array_obj_ref_343_final_offset) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_343_final_offset;
      ov(4 downto 0) := iv;
      array_obj_ref_343_root_address <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_addr_0
    process(array_obj_ref_349_root_address) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_349_root_address;
      ov(4 downto 0) := iv;
      array_obj_ref_349_word_address_0 <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_gather_scatter
    process(val_odd_341) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := val_odd_341;
      ov(31 downto 0) := iv;
      array_obj_ref_349_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_index_0_rename
    process(ADD_u8_u8_348_resized) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u8_u8_348_resized;
      ov(4 downto 0) := iv;
      ADD_u8_u8_348_scaled <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_index_0_resize
    process(ADD_u8_u8_348_wire) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u8_u8_348_wire;
      ov := iv(4 downto 0);
      ADD_u8_u8_348_resized <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_index_offset
    process(ADD_u8_u8_348_scaled) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u8_u8_348_scaled;
      ov(4 downto 0) := iv;
      array_obj_ref_349_final_offset <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_349_root_address_inst
    process(array_obj_ref_349_final_offset) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_349_final_offset;
      ov(4 downto 0) := iv;
      array_obj_ref_349_root_address <= ov(4 downto 0);
      --
    end process;
    if_stmt_357_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_360_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_357_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_357_branch_req_0,
          ack0 => if_stmt_357_branch_ack_0,
          ack1 => if_stmt_357_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u8_u8_339_inst
    process(R_328) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(R_328, konst_338_wire_constant, tmp_var);
      ADD_u8_u8_339_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_348_inst
    process(R_328) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(R_328, konst_347_wire_constant, tmp_var);
      ADD_u8_u8_348_wire <= tmp_var; --
    end process;
    -- shared split operator group (2) : ADD_u8_u8_355_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_328;
      nR_356 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_355_inst_req_0;
      ADD_u8_u8_355_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_355_inst_req_1;
      ADD_u8_u8_355_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator ULT_u8_u1_360_inst
    process(nR_356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nR_356, konst_359_wire_constant, tmp_var);
      ULT_u8_u1_360_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_349_store_0 array_obj_ref_343_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= array_obj_ref_349_store_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_343_store_0_req_0;
      array_obj_ref_349_store_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_343_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= array_obj_ref_349_store_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_343_store_0_req_1;
      array_obj_ref_349_store_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_343_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_349_word_address_0 & array_obj_ref_343_word_address_0;
      data_in <= array_obj_ref_349_data_0 & array_obj_ref_343_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 5,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(4 downto 0),
          mdata => memory_space_8_sr_data(31 downto 0),
          mtag => memory_space_8_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared call operator group (0) : call_stmt_336_call 
    dotP_even_call_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_336_call_req_0;
      call_stmt_336_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_336_call_req_1;
      call_stmt_336_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      dotP_even_call_group_0_gI: SplitGuardInterface generic map(name => "dotP_even_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_328;
      val_even_336 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 8,
        owidth => 8,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => dotP_even_call_reqs(0),
          ackR => dotP_even_call_acks(0),
          dataR => dotP_even_call_data(7 downto 0),
          tagR => dotP_even_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => dotP_even_return_acks(0), -- cross-over
          ackL => dotP_even_return_reqs(0), -- cross-over
          dataL => dotP_even_return_data(31 downto 0),
          tagL => dotP_even_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_341_call 
    dotP_odd_call_group_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_341_call_req_0;
      call_stmt_341_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_341_call_req_1;
      call_stmt_341_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      dotP_odd_call_group_1_gI: SplitGuardInterface generic map(name => "dotP_odd_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ADD_u8_u8_339_wire;
      val_odd_341 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 8,
        owidth => 8,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => dotP_odd_call_reqs(0),
          ackR => dotP_odd_call_acks(0),
          dataR => dotP_odd_call_data(7 downto 0),
          tagR => dotP_odd_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => dotP_odd_return_acks(0), -- cross-over
          ackL => dotP_odd_return_reqs(0), -- cross-over
          dataL => dotP_odd_return_data(31 downto 0),
          tagL => dotP_odd_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end multiplyMatrixVector_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity mvp_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    readVector_call_reqs : out  std_logic_vector(0 downto 0);
    readVector_call_acks : in   std_logic_vector(0 downto 0);
    readVector_call_tag  :  out  std_logic_vector(0 downto 0);
    readVector_return_reqs : out  std_logic_vector(0 downto 0);
    readVector_return_acks : in   std_logic_vector(0 downto 0);
    readVector_return_tag :  in   std_logic_vector(0 downto 0);
    multiplyMatrixVector_call_reqs : out  std_logic_vector(0 downto 0);
    multiplyMatrixVector_call_acks : in   std_logic_vector(0 downto 0);
    multiplyMatrixVector_call_tag  :  out  std_logic_vector(0 downto 0);
    multiplyMatrixVector_return_reqs : out  std_logic_vector(0 downto 0);
    multiplyMatrixVector_return_acks : in   std_logic_vector(0 downto 0);
    multiplyMatrixVector_return_tag :  in   std_logic_vector(0 downto 0);
    readMatrix_call_reqs : out  std_logic_vector(0 downto 0);
    readMatrix_call_acks : in   std_logic_vector(0 downto 0);
    readMatrix_call_tag  :  out  std_logic_vector(0 downto 0);
    readMatrix_return_reqs : out  std_logic_vector(0 downto 0);
    readMatrix_return_acks : in   std_logic_vector(0 downto 0);
    readMatrix_return_tag :  in   std_logic_vector(0 downto 0);
    sendVector_call_reqs : out  std_logic_vector(0 downto 0);
    sendVector_call_acks : in   std_logic_vector(0 downto 0);
    sendVector_call_tag  :  out  std_logic_vector(0 downto 0);
    sendVector_return_reqs : out  std_logic_vector(0 downto 0);
    sendVector_return_acks : in   std_logic_vector(0 downto 0);
    sendVector_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mvp_daemon;
architecture mvp_daemon_arch of mvp_daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal mvp_daemon_CP_3398_start: Boolean;
  signal mvp_daemon_CP_3398_symbol: Boolean;
  -- volatile/operator module components. 
  component readVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component multiplyMatrixVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      dotP_even_call_reqs : out  std_logic_vector(0 downto 0);
      dotP_even_call_acks : in   std_logic_vector(0 downto 0);
      dotP_even_call_data : out  std_logic_vector(7 downto 0);
      dotP_even_call_tag  :  out  std_logic_vector(0 downto 0);
      dotP_even_return_reqs : out  std_logic_vector(0 downto 0);
      dotP_even_return_acks : in   std_logic_vector(0 downto 0);
      dotP_even_return_data : in   std_logic_vector(31 downto 0);
      dotP_even_return_tag :  in   std_logic_vector(0 downto 0);
      dotP_odd_call_reqs : out  std_logic_vector(0 downto 0);
      dotP_odd_call_acks : in   std_logic_vector(0 downto 0);
      dotP_odd_call_data : out  std_logic_vector(7 downto 0);
      dotP_odd_call_tag  :  out  std_logic_vector(0 downto 0);
      dotP_odd_return_reqs : out  std_logic_vector(0 downto 0);
      dotP_odd_return_acks : in   std_logic_vector(0 downto 0);
      dotP_odd_return_data : in   std_logic_vector(31 downto 0);
      dotP_odd_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component readMatrix is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(4 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_610_call_ack_0 : boolean;
  signal call_stmt_612_call_req_0 : boolean;
  signal call_stmt_610_call_ack_1 : boolean;
  signal call_stmt_607_call_req_1 : boolean;
  signal call_stmt_610_call_req_0 : boolean;
  signal call_stmt_607_call_ack_1 : boolean;
  signal call_stmt_610_call_req_1 : boolean;
  signal call_stmt_612_call_ack_0 : boolean;
  signal call_stmt_612_call_ack_1 : boolean;
  signal call_stmt_612_call_req_1 : boolean;
  signal call_stmt_611_call_req_0 : boolean;
  signal call_stmt_607_call_ack_0 : boolean;
  signal call_stmt_611_call_ack_1 : boolean;
  signal call_stmt_611_call_req_1 : boolean;
  signal call_stmt_607_call_req_0 : boolean;
  signal call_stmt_611_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "mvp_daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  mvp_daemon_CP_3398_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "mvp_daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mvp_daemon_CP_3398_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= mvp_daemon_CP_3398_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mvp_daemon_CP_3398_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  mvp_daemon_CP_3398: Block -- control-path 
    signal mvp_daemon_CP_3398_elements: BooleanArray(12 downto 0);
    -- 
  begin -- 
    mvp_daemon_CP_3398_elements(0) <= mvp_daemon_CP_3398_start;
    mvp_daemon_CP_3398_symbol <= mvp_daemon_CP_3398_elements(3);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_Update/ccr
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_Sample/$entry
      -- CP-element group 0: 	 call_stmt_607/$entry
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_sample_start_
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_update_start_
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_Update/$entry
      -- CP-element group 0: 	 call_stmt_607/call_stmt_607_Sample/crr
      -- 
    crr_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(0), ack => call_stmt_607_call_req_0); -- 
    ccr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(0), ack => call_stmt_607_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_607/call_stmt_607_sample_completed_
      -- CP-element group 1: 	 call_stmt_607/call_stmt_607_Sample/cra
      -- CP-element group 1: 	 call_stmt_607/call_stmt_607_Sample/$exit
      -- 
    cra_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_607_call_ack_0, ack => mvp_daemon_CP_3398_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_608/branch_block_stmt_608__entry__
      -- CP-element group 2: 	 call_stmt_607/call_stmt_607_update_completed_
      -- CP-element group 2: 	 call_stmt_607/call_stmt_607_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_608/merge_stmt_609__entry__
      -- CP-element group 2: 	 branch_block_stmt_608/$entry
      -- CP-element group 2: 	 call_stmt_607/$exit
      -- CP-element group 2: 	 call_stmt_607/call_stmt_607_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_608/merge_stmt_609__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_608/merge_stmt_609__entry___PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_608/merge_stmt_609_dead_link/$entry
      -- 
    cca_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_607_call_ack_1, ack => mvp_daemon_CP_3398_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_608/$exit
      -- CP-element group 3: 	 branch_block_stmt_608/branch_block_stmt_608__exit__
      -- 
    mvp_daemon_CP_3398_elements(3) <= false; 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	12 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Sample/cra
      -- CP-element group 4: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_sample_completed_
      -- 
    cra_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_610_call_ack_0, ack => mvp_daemon_CP_3398_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	12 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	10 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Update/cca
      -- CP-element group 5: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_update_completed_
      -- 
    cca_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_610_call_ack_1, ack => mvp_daemon_CP_3398_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	10 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Sample/cra
      -- 
    cra_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_611_call_ack_0, ack => mvp_daemon_CP_3398_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	11 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Update/cca
      -- CP-element group 7: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Update/$exit
      -- 
    cca_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_611_call_ack_1, ack => mvp_daemon_CP_3398_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Sample/cra
      -- CP-element group 8: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_sample_completed_
      -- 
    cra_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_612_call_ack_0, ack => mvp_daemon_CP_3398_elements(8)); -- 
    -- CP-element group 9:  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (8) 
      -- CP-element group 9: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/$exit
      -- CP-element group 9: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612__exit__
      -- CP-element group 9: 	 branch_block_stmt_608/loopback
      -- CP-element group 9: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Update/cca
      -- CP-element group 9: 	 branch_block_stmt_608/loopback_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_608/loopback_PhiReq/$exit
      -- 
    cca_3472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_612_call_ack_1, ack => mvp_daemon_CP_3398_elements(9)); -- 
    -- CP-element group 10:  transition  output  delay-element  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	5 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	6 
    -- CP-element group 10:  members (4) 
      -- CP-element group 10: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Sample/crr
      -- CP-element group 10: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_call_stmt_611_delay
      -- 
    crr_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(10), ack => call_stmt_611_call_req_0); -- 
    -- Element group mvp_daemon_CP_3398_elements(10) is a control-delay.
    cp_element_10_delay: control_delay_element  generic map(name => " 10_delay", delay_value => 1)  port map(req => mvp_daemon_CP_3398_elements(5), ack => mvp_daemon_CP_3398_elements(10), clk => clk, reset =>reset);
    -- CP-element group 11:  transition  output  delay-element  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	7 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	8 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Sample/crr
      -- CP-element group 11: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_call_stmt_612_delay
      -- 
    crr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(11), ack => call_stmt_612_call_req_0); -- 
    -- Element group mvp_daemon_CP_3398_elements(11) is a control-delay.
    cp_element_11_delay: control_delay_element  generic map(name => " 11_delay", delay_value => 1)  port map(req => mvp_daemon_CP_3398_elements(7), ack => mvp_daemon_CP_3398_elements(11), clk => clk, reset =>reset);
    -- CP-element group 12:  merge  fork  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	5 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	4 
    -- CP-element group 12: 	9 
    -- CP-element group 12:  members (19) 
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/merge_stmt_609__exit__
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612__entry__
      -- CP-element group 12: 	 branch_block_stmt_608/merge_stmt_609_PhiReqMerge
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_update_start_
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_update_start_
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Sample/crr
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_Update/ccr
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_612_Update/ccr
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_610_update_start_
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Update/ccr
      -- CP-element group 12: 	 branch_block_stmt_608/call_stmt_610_to_call_stmt_612/call_stmt_611_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/merge_stmt_609_PhiAck/dummy
      -- CP-element group 12: 	 branch_block_stmt_608/merge_stmt_609_PhiAck/$entry
      -- CP-element group 12: 	 branch_block_stmt_608/merge_stmt_609_PhiAck/$exit
      -- 
    crr_3438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(12), ack => call_stmt_610_call_req_0); -- 
    ccr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(12), ack => call_stmt_610_call_req_1); -- 
    ccr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(12), ack => call_stmt_612_call_req_1); -- 
    ccr_3457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mvp_daemon_CP_3398_elements(12), ack => call_stmt_611_call_req_1); -- 
    mvp_daemon_CP_3398_elements(12) <= OrReduce(mvp_daemon_CP_3398_elements(9) & mvp_daemon_CP_3398_elements(2));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_607_call 
    readMatrix_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_607_call_req_0;
      call_stmt_607_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_607_call_req_1;
      call_stmt_607_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readMatrix_call_group_0_gI: SplitGuardInterface generic map(name => "readMatrix_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => readMatrix_call_reqs(0),
          ackR => readMatrix_call_acks(0),
          tagR => readMatrix_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => readMatrix_return_acks(0), -- cross-over
          ackL => readMatrix_return_reqs(0), -- cross-over
          tagL => readMatrix_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_610_call 
    readVector_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_610_call_req_0;
      call_stmt_610_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_610_call_req_1;
      call_stmt_610_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readVector_call_group_1_gI: SplitGuardInterface generic map(name => "readVector_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => readVector_call_reqs(0),
          ackR => readVector_call_acks(0),
          tagR => readVector_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => readVector_return_acks(0), -- cross-over
          ackL => readVector_return_reqs(0), -- cross-over
          tagL => readVector_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_611_call 
    multiplyMatrixVector_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_611_call_req_0;
      call_stmt_611_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_611_call_req_1;
      call_stmt_611_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      multiplyMatrixVector_call_group_2_gI: SplitGuardInterface generic map(name => "multiplyMatrixVector_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => multiplyMatrixVector_call_reqs(0),
          ackR => multiplyMatrixVector_call_acks(0),
          tagR => multiplyMatrixVector_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => multiplyMatrixVector_return_acks(0), -- cross-over
          ackL => multiplyMatrixVector_return_reqs(0), -- cross-over
          tagL => multiplyMatrixVector_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_612_call 
    sendVector_call_group_3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_612_call_req_0;
      call_stmt_612_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_612_call_req_1;
      call_stmt_612_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendVector_call_group_3_gI: SplitGuardInterface generic map(name => "sendVector_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendVector_call_reqs(0),
          ackR => sendVector_call_acks(0),
          tagR => sendVector_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendVector_return_acks(0), -- cross-over
          ackL => sendVector_return_reqs(0), -- cross-over
          tagL => sendVector_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end mvp_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readMatrix is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readMatrix;
architecture readMatrix_arch of readMatrix is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal readMatrix_CP_2257_start: Boolean;
  signal readMatrix_CP_2257_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_450_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_426_store_0_ack_0 : boolean;
  signal array_obj_ref_426_store_0_req_0 : boolean;
  signal slice_398_inst_req_1 : boolean;
  signal array_obj_ref_450_index_0_scale_req_0 : boolean;
  signal array_obj_ref_450_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_450_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_450_index_sum_1_req_1 : boolean;
  signal ADD_u8_u8_377_inst_ack_0 : boolean;
  signal array_obj_ref_438_index_0_scale_ack_0 : boolean;
  signal ADD_u8_u8_377_inst_req_0 : boolean;
  signal array_obj_ref_426_index_sum_1_req_0 : boolean;
  signal array_obj_ref_438_index_sum_1_req_1 : boolean;
  signal array_obj_ref_426_index_sum_1_ack_1 : boolean;
  signal RPIPE_in_data_401_inst_req_0 : boolean;
  signal array_obj_ref_450_store_0_req_0 : boolean;
  signal array_obj_ref_450_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_450_index_sum_1_req_0 : boolean;
  signal array_obj_ref_438_index_0_scale_req_0 : boolean;
  signal array_obj_ref_450_store_0_ack_0 : boolean;
  signal array_obj_ref_438_store_0_ack_1 : boolean;
  signal array_obj_ref_426_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_426_index_0_scale_req_1 : boolean;
  signal array_obj_ref_426_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_426_index_sum_1_req_1 : boolean;
  signal array_obj_ref_426_index_0_scale_req_0 : boolean;
  signal array_obj_ref_450_store_0_req_1 : boolean;
  signal array_obj_ref_462_index_0_scale_req_1 : boolean;
  signal array_obj_ref_438_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_1 : boolean;
  signal RPIPE_in_data_401_inst_ack_0 : boolean;
  signal slice_398_inst_ack_0 : boolean;
  signal array_obj_ref_438_index_sum_1_req_0 : boolean;
  signal array_obj_ref_462_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_438_store_0_req_0 : boolean;
  signal array_obj_ref_462_index_0_scale_req_0 : boolean;
  signal array_obj_ref_438_index_sum_1_ack_1 : boolean;
  signal ADD_u8_u8_377_inst_req_1 : boolean;
  signal array_obj_ref_462_index_0_scale_ack_0 : boolean;
  signal ADD_u8_u8_377_inst_ack_1 : boolean;
  signal array_obj_ref_450_index_0_scale_req_1 : boolean;
  signal array_obj_ref_450_store_0_ack_1 : boolean;
  signal array_obj_ref_426_index_sum_1_ack_0 : boolean;
  signal slice_398_inst_ack_1 : boolean;
  signal array_obj_ref_438_store_0_ack_0 : boolean;
  signal ADD_u8_u8_389_inst_ack_1 : boolean;
  signal ADD_u8_u8_389_inst_req_1 : boolean;
  signal ADD_u8_u8_389_inst_ack_0 : boolean;
  signal ADD_u8_u8_389_inst_req_0 : boolean;
  signal array_obj_ref_426_store_0_ack_1 : boolean;
  signal slice_398_inst_req_0 : boolean;
  signal array_obj_ref_426_store_0_req_1 : boolean;
  signal array_obj_ref_438_index_0_scale_ack_1 : boolean;
  signal RPIPE_in_data_401_inst_ack_1 : boolean;
  signal RPIPE_in_data_401_inst_req_1 : boolean;
  signal array_obj_ref_438_index_0_scale_req_1 : boolean;
  signal array_obj_ref_462_index_sum_1_req_0 : boolean;
  signal array_obj_ref_462_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_462_index_sum_1_req_1 : boolean;
  signal array_obj_ref_462_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_462_store_0_req_0 : boolean;
  signal array_obj_ref_462_store_0_ack_0 : boolean;
  signal array_obj_ref_462_store_0_req_1 : boolean;
  signal array_obj_ref_462_store_0_ack_1 : boolean;
  signal if_stmt_471_branch_req_0 : boolean;
  signal if_stmt_471_branch_ack_1 : boolean;
  signal if_stmt_471_branch_ack_0 : boolean;
  signal if_stmt_477_branch_req_0 : boolean;
  signal if_stmt_477_branch_ack_1 : boolean;
  signal if_stmt_477_branch_ack_0 : boolean;
  signal phi_stmt_368_req_0 : boolean;
  signal nI_378_372_buf_req_0 : boolean;
  signal nI_378_372_buf_ack_0 : boolean;
  signal nI_378_372_buf_req_1 : boolean;
  signal nI_378_372_buf_ack_1 : boolean;
  signal phi_stmt_368_req_1 : boolean;
  signal phi_stmt_368_ack_0 : boolean;
  signal phi_stmt_380_req_0 : boolean;
  signal nJ_390_384_buf_req_0 : boolean;
  signal nJ_390_384_buf_ack_0 : boolean;
  signal nJ_390_384_buf_req_1 : boolean;
  signal nJ_390_384_buf_ack_1 : boolean;
  signal phi_stmt_380_req_1 : boolean;
  signal phi_stmt_380_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readMatrix_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readMatrix_CP_2257_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readMatrix_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readMatrix_CP_2257_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readMatrix_CP_2257_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readMatrix_CP_2257_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readMatrix_CP_2257: Block -- control-path 
    signal readMatrix_CP_2257_elements: BooleanArray(57 downto 0);
    -- 
  begin -- 
    readMatrix_CP_2257_elements(0) <= readMatrix_CP_2257_start;
    readMatrix_CP_2257_symbol <= readMatrix_CP_2257_elements(45);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	46 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_366/$entry
      -- CP-element group 0: 	 branch_block_stmt_366/merge_stmt_367__entry__
      -- CP-element group 0: 	 branch_block_stmt_366/branch_block_stmt_366__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_366/merge_stmt_367_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/$entry
      -- CP-element group 0: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/phi_stmt_368_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	51 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_sample_completed_
      -- 
    ra_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_377_inst_ack_0, ack => readMatrix_CP_2257_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	51 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	52 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_366/merge_stmt_379__entry__
      -- CP-element group 2: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_366/assign_stmt_378/$exit
      -- CP-element group 2: 	 branch_block_stmt_366/assign_stmt_378__exit__
      -- CP-element group 2: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_366/merge_stmt_379_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/$entry
      -- CP-element group 2: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/phi_stmt_380_sources/$entry
      -- 
    ca_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_377_inst_ack_1, ack => readMatrix_CP_2257_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	57 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_sample_completed_
      -- 
    ra_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_389_inst_ack_0, ack => readMatrix_CP_2257_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	57 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	41 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_update_completed_
      -- 
    ca_2310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u8_u8_389_inst_ack_1, ack => readMatrix_CP_2257_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	57 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_sample_completed_
      -- 
    ra_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_398_inst_ack_0, ack => readMatrix_CP_2257_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	57 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	12 
    -- CP-element group 6: 	20 
    -- CP-element group 6: 	28 
    -- CP-element group 6: 	36 
    -- CP-element group 6:  members (47) 
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scaled_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_1/index_resize_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scaled_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resized_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_computed_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resized_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scaled_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resized_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_computed_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_1/index_resize_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_computed_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scaled_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resized_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_1/index_resize_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_1/$exit
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_computed_1
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_1/index_resize_req
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_1/$entry
      -- CP-element group 6: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_1/$exit
      -- 
    ca_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_398_inst_ack_1, ack => readMatrix_CP_2257_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	57 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_update_start_
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Update/cr
      -- 
    ra_2333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_401_inst_ack_0, ack => readMatrix_CP_2257_elements(7)); -- 
    cr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(7), ack => RPIPE_in_data_401_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	33 
    -- CP-element group 8: 	25 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Update/ca
      -- 
    ca_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_401_inst_ack_1, ack => readMatrix_CP_2257_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/word_0/rr
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/array_obj_ref_426_Split/split_ack
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/array_obj_ref_426_Split/split_req
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/word_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/$entry
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/array_obj_ref_426_Split/$exit
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/array_obj_ref_426_Split/$entry
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_sample_start_
      -- 
    rr_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(9), ack => array_obj_ref_426_store_0_req_0); -- 
    readMatrix_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "readMatrix_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(14) & readMatrix_CP_2257_elements(8);
      gj_readMatrix_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	57 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	41 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_sample_complete
      -- 
    ra_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_index_0_scale_ack_0, ack => readMatrix_CP_2257_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	57 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (4) 
      -- CP-element group 11: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_update_complete
      -- CP-element group 11: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scaled_0
      -- 
    ca_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_index_0_scale_ack_1, ack => readMatrix_CP_2257_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: 	6 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_sample_start
      -- 
    rr_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(12), ack => array_obj_ref_426_index_sum_1_req_0); -- 
    readMatrix_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(11) & readMatrix_CP_2257_elements(6);
      gj_readMatrix_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_sample_complete
      -- CP-element group 13: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Sample/ra
      -- 
    ra_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_index_sum_1_ack_0, ack => readMatrix_CP_2257_elements(13)); -- 
    -- CP-element group 14:  join  fork  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	57 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (18) 
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_update_complete
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_final_index_sum_regn/$entry
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_word_addrgen/root_register_ack
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_word_addrgen/root_register_req
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_word_addrgen/$exit
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_word_addrgen/$entry
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_offset_calculated
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_root_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_word_address_calculated
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_base_plus_offset/$exit
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_base_plus_offset/$entry
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_final_index_sum_regn/ack
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_final_index_sum_regn/req
      -- CP-element group 14: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_final_index_sum_regn/$exit
      -- 
    ca_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_index_sum_1_ack_1, ack => readMatrix_CP_2257_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_sample_completed_
      -- 
    ra_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_store_0_ack_0, ack => readMatrix_CP_2257_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/$exit
      -- 
    ca_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_426_store_0_ack_1, ack => readMatrix_CP_2257_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	22 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/array_obj_ref_438_Split/split_req
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/array_obj_ref_438_Split/$exit
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/array_obj_ref_438_Split/split_ack
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/word_0/rr
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/array_obj_ref_438_Split/$entry
      -- CP-element group 17: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_sample_start_
      -- 
    rr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(17), ack => array_obj_ref_438_store_0_req_0); -- 
    readMatrix_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(8) & readMatrix_CP_2257_elements(22);
      gj_readMatrix_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	57 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_sample_complete
      -- 
    ra_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_index_0_scale_ack_0, ack => readMatrix_CP_2257_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	57 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_update_complete
      -- CP-element group 19: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scaled_0
      -- CP-element group 19: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Update/$exit
      -- 
    ca_2465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_index_0_scale_ack_1, ack => readMatrix_CP_2257_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_sample_start
      -- 
    rr_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(20), ack => array_obj_ref_438_index_sum_1_req_0); -- 
    readMatrix_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(6) & readMatrix_CP_2257_elements(19);
      gj_readMatrix_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_sample_complete
      -- 
    ra_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_index_sum_1_ack_0, ack => readMatrix_CP_2257_elements(21)); -- 
    -- CP-element group 22:  join  fork  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	57 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (18) 
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_base_plus_offset/$exit
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_final_index_sum_regn/ack
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_word_addrgen/$exit
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_word_addrgen/root_register_req
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_base_plus_offset/$entry
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_final_index_sum_regn/$entry
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_final_index_sum_regn/req
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_final_index_sum_regn/$exit
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_root_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_offset_calculated
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_update_complete
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_word_address_calculated
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_word_addrgen/$entry
      -- CP-element group 22: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_word_addrgen/root_register_ack
      -- 
    ca_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_index_sum_1_ack_1, ack => readMatrix_CP_2257_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_sample_completed_
      -- 
    ra_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_0, ack => readMatrix_CP_2257_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	57 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	41 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/$exit
      -- 
    ca_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_1, ack => readMatrix_CP_2257_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	8 
    -- CP-element group 25: 	30 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/word_0/rr
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/array_obj_ref_450_Split/$exit
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/array_obj_ref_450_Split/$entry
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/word_0/$entry
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/array_obj_ref_450_Split/split_req
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/array_obj_ref_450_Split/split_ack
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/$entry
      -- CP-element group 25: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/$entry
      -- 
    rr_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(25), ack => array_obj_ref_450_store_0_req_0); -- 
    readMatrix_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(8) & readMatrix_CP_2257_elements(30);
      gj_readMatrix_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	57 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	41 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_sample_complete
      -- CP-element group 26: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Sample/$exit
      -- 
    ra_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_index_0_scale_ack_0, ack => readMatrix_CP_2257_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	57 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_update_complete
      -- CP-element group 27: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scaled_0
      -- 
    ca_2563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_index_0_scale_ack_1, ack => readMatrix_CP_2257_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	6 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_sample_start
      -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(28), ack => array_obj_ref_450_index_sum_1_req_0); -- 
    readMatrix_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(6) & readMatrix_CP_2257_elements(27);
      gj_readMatrix_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	41 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_sample_complete
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_index_sum_1_ack_0, ack => readMatrix_CP_2257_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	57 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	25 
    -- CP-element group 30:  members (18) 
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_root_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_base_plus_offset/$entry
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_final_index_sum_regn/$exit
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_base_plus_offset/$exit
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_final_index_sum_regn/$entry
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_word_addrgen/$entry
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_update_complete
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_word_address_calculated
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_final_index_sum_regn/ack
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_final_index_sum_regn/req
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_word_addrgen/root_register_ack
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_word_addrgen/root_register_req
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_offset_calculated
      -- CP-element group 30: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_word_addrgen/$exit
      -- 
    ca_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_index_sum_1_ack_1, ack => readMatrix_CP_2257_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	25 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/word_0/ra
      -- CP-element group 31: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Sample/$exit
      -- 
    ra_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_store_0_ack_0, ack => readMatrix_CP_2257_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	41 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/word_0/ca
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_store_0_ack_1, ack => readMatrix_CP_2257_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	8 
    -- CP-element group 33: 	38 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	39 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/array_obj_ref_462_Split/$entry
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/array_obj_ref_462_Split/$exit
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/array_obj_ref_462_Split/split_req
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/array_obj_ref_462_Split/split_ack
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/word_0/rr
      -- 
    rr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(33), ack => array_obj_ref_462_store_0_req_0); -- 
    readMatrix_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(8) & readMatrix_CP_2257_elements(38);
      gj_readMatrix_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	57 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_sample_complete
      -- CP-element group 34: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Sample/ra
      -- 
    ra_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_0_scale_ack_0, ack => readMatrix_CP_2257_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	57 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_update_complete
      -- CP-element group 35: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scaled_0
      -- 
    ca_2661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_0_scale_ack_1, ack => readMatrix_CP_2257_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	6 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_sample_start
      -- CP-element group 36: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Sample/$entry
      -- 
    rr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(36), ack => array_obj_ref_462_index_sum_1_req_0); -- 
    readMatrix_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(6) & readMatrix_CP_2257_elements(35);
      gj_readMatrix_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	41 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_sample_complete
      -- CP-element group 37: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Sample/$exit
      -- 
    ra_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_sum_1_ack_0, ack => readMatrix_CP_2257_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	33 
    -- CP-element group 38:  members (18) 
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_offset_calculated
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_word_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_root_address_calculated
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_base_plus_offset/sum_rename_req
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_base_plus_offset/sum_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_base_plus_offset/$entry
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_base_plus_offset/$exit
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_final_index_sum_regn/$entry
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_final_index_sum_regn/req
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_final_index_sum_regn/ack
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_final_index_sum_regn/$exit
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_update_complete
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_word_addrgen/$entry
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_word_addrgen/$exit
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_word_addrgen/root_register_req
      -- CP-element group 38: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_word_addrgen/root_register_ack
      -- 
    ca_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_sum_1_ack_1, ack => readMatrix_CP_2257_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	33 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/$exit
      -- CP-element group 39: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Sample/word_access_start/word_0/ra
      -- 
    ra_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_store_0_ack_0, ack => readMatrix_CP_2257_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	57 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/$exit
      -- CP-element group 40: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/word_0/ca
      -- 
    ca_2730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_store_0_ack_1, ack => readMatrix_CP_2257_elements(40)); -- 
    -- CP-element group 41:  branch  join  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: 	10 
    -- CP-element group 41: 	4 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	32 
    -- CP-element group 41: 	34 
    -- CP-element group 41: 	29 
    -- CP-element group 41: 	26 
    -- CP-element group 41: 	24 
    -- CP-element group 41: 	37 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (24) 
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471__entry__
      -- CP-element group 41: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464__exit__
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_dead_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/ULT_u8_u1_474_inputs/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/ULT_u8_u1_474_inputs/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Update/cr
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/ULT_u8_u1_474/SplitProtocol/Update/ca
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_eval_test/branch_req
      -- CP-element group 41: 	 branch_block_stmt_366/ULT_u8_u1_474_place
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_if_link/$entry
      -- CP-element group 41: 	 branch_block_stmt_366/if_stmt_471_else_link/$entry
      -- 
    branch_req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(41), ack => if_stmt_471_branch_req_0); -- 
    readMatrix_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(13) & readMatrix_CP_2257_elements(10) & readMatrix_CP_2257_elements(4) & readMatrix_CP_2257_elements(16) & readMatrix_CP_2257_elements(18) & readMatrix_CP_2257_elements(21) & readMatrix_CP_2257_elements(32) & readMatrix_CP_2257_elements(34) & readMatrix_CP_2257_elements(29) & readMatrix_CP_2257_elements(26) & readMatrix_CP_2257_elements(24) & readMatrix_CP_2257_elements(37) & readMatrix_CP_2257_elements(40);
      gj_readMatrix_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  place  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	53 
    -- CP-element group 42: 	54 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_366/if_stmt_471_if_link/$exit
      -- CP-element group 42: 	 branch_block_stmt_366/if_stmt_471_if_link/if_choice_transition
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Sample/req
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Update/req
      -- 
    if_choice_transition_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_471_branch_ack_1, ack => readMatrix_CP_2257_elements(42)); -- 
    req_2878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(42), ack => nJ_390_384_buf_req_0); -- 
    req_2883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(42), ack => nJ_390_384_buf_req_1); -- 
    -- CP-element group 43:  merge  branch  transition  place  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (25) 
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477__entry__
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_471__exit__
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_471_else_link/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_471_else_link/else_choice_transition
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_dead_link/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/ULT_u8_u1_480_inputs/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/ULT_u8_u1_480_inputs/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/ULT_u8_u1_480/SplitProtocol/Update/ca
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_eval_test/branch_req
      -- CP-element group 43: 	 branch_block_stmt_366/ULT_u8_u1_480_place
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_if_link/$entry
      -- CP-element group 43: 	 branch_block_stmt_366/if_stmt_477_else_link/$entry
      -- 
    else_choice_transition_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_471_branch_ack_0, ack => readMatrix_CP_2257_elements(43)); -- 
    branch_req_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(43), ack => if_stmt_477_branch_req_0); -- 
    -- CP-element group 44:  fork  transition  place  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: 	48 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_366/if_stmt_477_if_link/$exit
      -- CP-element group 44: 	 branch_block_stmt_366/if_stmt_477_if_link/if_choice_transition
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Sample/req
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Update/req
      -- 
    if_choice_transition_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_477_branch_ack_1, ack => readMatrix_CP_2257_elements(44)); -- 
    req_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(44), ack => nI_378_372_buf_req_0); -- 
    req_2840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(44), ack => nI_378_372_buf_req_1); -- 
    -- CP-element group 45:  merge  transition  place  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_366/if_stmt_477__exit__
      -- CP-element group 45: 	 $exit
      -- CP-element group 45: 	 branch_block_stmt_366/$exit
      -- CP-element group 45: 	 branch_block_stmt_366/branch_block_stmt_366__exit__
      -- CP-element group 45: 	 branch_block_stmt_366/if_stmt_477_else_link/$exit
      -- CP-element group 45: 	 branch_block_stmt_366/if_stmt_477_else_link/else_choice_transition
      -- 
    else_choice_transition_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_477_branch_ack_0, ack => readMatrix_CP_2257_elements(45)); -- 
    -- CP-element group 46:  transition  output  delay-element  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	0 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	50 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/$exit
      -- CP-element group 46: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/$exit
      -- CP-element group 46: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/phi_stmt_368_sources/$exit
      -- CP-element group 46: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/phi_stmt_368_sources/type_cast_371_konst_delay_trans
      -- CP-element group 46: 	 branch_block_stmt_366/merge_stmt_367__entry___PhiReq/phi_stmt_368/phi_stmt_368_req
      -- 
    phi_stmt_368_req_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_368_req_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(46), ack => phi_stmt_368_req_0); -- 
    -- Element group readMatrix_CP_2257_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => readMatrix_CP_2257_elements(0), ack => readMatrix_CP_2257_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Sample/ack
      -- 
    ack_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_378_372_buf_ack_0, ack => readMatrix_CP_2257_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	44 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/Update/ack
      -- 
    ack_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_378_372_buf_ack_1, ack => readMatrix_CP_2257_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_366/outer_loopback_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/$exit
      -- CP-element group 49: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/$exit
      -- CP-element group 49: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_sources/Interlock/$exit
      -- CP-element group 49: 	 branch_block_stmt_366/outer_loopback_PhiReq/phi_stmt_368/phi_stmt_368_req
      -- 
    phi_stmt_368_req_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_368_req_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(49), ack => phi_stmt_368_req_1); -- 
    readMatrix_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(47) & readMatrix_CP_2257_elements(48);
      gj_readMatrix_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  merge  transition  place  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	46 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_366/merge_stmt_367_PhiReqMerge
      -- CP-element group 50: 	 branch_block_stmt_366/merge_stmt_367_PhiAck/$entry
      -- 
    readMatrix_CP_2257_elements(50) <= OrReduce(readMatrix_CP_2257_elements(46) & readMatrix_CP_2257_elements(49));
    -- CP-element group 51:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	1 
    -- CP-element group 51: 	2 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/$entry
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_update_start_
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378__entry__
      -- CP-element group 51: 	 branch_block_stmt_366/merge_stmt_367__exit__
      -- CP-element group 51: 	 branch_block_stmt_366/assign_stmt_378/ADD_u8_u8_377_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_366/merge_stmt_367_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_366/merge_stmt_367_PhiAck/phi_stmt_368_ack
      -- 
    phi_stmt_368_ack_2847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_368_ack_0, ack => readMatrix_CP_2257_elements(51)); -- 
    rr_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(51), ack => ADD_u8_u8_377_inst_req_0); -- 
    cr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(51), ack => ADD_u8_u8_377_inst_req_1); -- 
    -- CP-element group 52:  transition  output  delay-element  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	2 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	56 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/$exit
      -- CP-element group 52: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/phi_stmt_380_sources/$exit
      -- CP-element group 52: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/phi_stmt_380_sources/type_cast_383_konst_delay_trans
      -- CP-element group 52: 	 branch_block_stmt_366/merge_stmt_379__entry___PhiReq/phi_stmt_380/phi_stmt_380_req
      -- 
    phi_stmt_380_req_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_380_req_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(52), ack => phi_stmt_380_req_0); -- 
    -- Element group readMatrix_CP_2257_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => readMatrix_CP_2257_elements(2), ack => readMatrix_CP_2257_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	42 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Sample/ack
      -- 
    ack_2879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nJ_390_384_buf_ack_0, ack => readMatrix_CP_2257_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	42 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/Update/ack
      -- 
    ack_2884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nJ_390_384_buf_ack_1, ack => readMatrix_CP_2257_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_366/inner_loopback_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/$exit
      -- CP-element group 55: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/$exit
      -- CP-element group 55: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_sources/Interlock/$exit
      -- CP-element group 55: 	 branch_block_stmt_366/inner_loopback_PhiReq/phi_stmt_380/phi_stmt_380_req
      -- 
    phi_stmt_380_req_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_380_req_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(55), ack => phi_stmt_380_req_1); -- 
    readMatrix_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readMatrix_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMatrix_CP_2257_elements(53) & readMatrix_CP_2257_elements(54);
      gj_readMatrix_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMatrix_CP_2257_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  transition  place  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_366/merge_stmt_379_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_366/merge_stmt_379_PhiAck/$entry
      -- 
    readMatrix_CP_2257_elements(56) <= OrReduce(readMatrix_CP_2257_elements(52) & readMatrix_CP_2257_elements(55));
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	3 
    -- CP-element group 57: 	11 
    -- CP-element group 57: 	14 
    -- CP-element group 57: 	10 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	5 
    -- CP-element group 57: 	6 
    -- CP-element group 57: 	7 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	18 
    -- CP-element group 57: 	19 
    -- CP-element group 57: 	22 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	34 
    -- CP-element group 57: 	30 
    -- CP-element group 57: 	26 
    -- CP-element group 57: 	27 
    -- CP-element group 57: 	24 
    -- CP-element group 57: 	35 
    -- CP-element group 57: 	38 
    -- CP-element group 57: 	40 
    -- CP-element group 57:  members (100) 
      -- CP-element group 57: 	 branch_block_stmt_366/merge_stmt_379__exit__
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464__entry__
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_sample_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_0/index_resize_ack
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_0/index_resize_req
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resize_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/word_0/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_0/index_resize_req
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_0/index_resize_ack
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/word_0/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resized_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_sample_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_sample_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_resized_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_partial_sum_1_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_0/index_resize_req
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_0/index_resize_ack
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_partial_sum_1_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_sample_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_0/index_resize_ack
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_scale_0_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_scale_0_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_0/index_resize_req
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_computed_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_scale_0_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_partial_sum_1_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resize_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_computed_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_index_resized_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resize_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/slice_398_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_computed_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/word_0/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/ADD_u8_u8_389_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_update_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/RPIPE_in_data_401_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_426_Update/word_access_complete/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_Update/word_access_complete/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_index_resized_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_438_index_scale_0_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_450_Update/word_access_complete/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_resize_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_update_start
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_index_computed_0
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_partial_sum_1_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/word_0/$entry
      -- CP-element group 57: 	 branch_block_stmt_366/assign_stmt_390_to_assign_stmt_464/array_obj_ref_462_Update/word_access_complete/word_0/cr
      -- CP-element group 57: 	 branch_block_stmt_366/merge_stmt_379_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_366/merge_stmt_379_PhiAck/phi_stmt_380_ack
      -- 
    phi_stmt_380_ack_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_380_ack_0, ack => readMatrix_CP_2257_elements(57)); -- 
    cr_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => slice_398_inst_req_1); -- 
    rr_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_450_index_0_scale_req_0); -- 
    cr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_450_index_sum_1_req_1); -- 
    cr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_438_index_sum_1_req_1); -- 
    rr_2332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => RPIPE_in_data_401_inst_req_0); -- 
    rr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_438_index_0_scale_req_0); -- 
    cr_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_426_index_0_scale_req_1); -- 
    cr_2393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_426_index_sum_1_req_1); -- 
    rr_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_426_index_0_scale_req_0); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_450_store_0_req_1); -- 
    cr_2660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_462_index_0_scale_req_1); -- 
    cr_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_438_store_0_req_1); -- 
    rr_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_462_index_0_scale_req_0); -- 
    cr_2562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_450_index_0_scale_req_1); -- 
    cr_2309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => ADD_u8_u8_389_inst_req_1); -- 
    rr_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => ADD_u8_u8_389_inst_req_0); -- 
    rr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => slice_398_inst_req_0); -- 
    cr_2435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_426_store_0_req_1); -- 
    cr_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_438_index_0_scale_req_1); -- 
    cr_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_462_index_sum_1_req_1); -- 
    cr_2729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMatrix_CP_2257_elements(57), ack => array_obj_ref_462_store_0_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_368 : std_logic_vector(7 downto 0);
    signal J_380 : std_logic_vector(7 downto 0);
    signal J_idx_0_407 : std_logic_vector(0 downto 0);
    signal J_idx_1_412 : std_logic_vector(0 downto 0);
    signal J_idx_2_417 : std_logic_vector(0 downto 0);
    signal J_idx_395 : std_logic_vector(1 downto 0);
    signal J_idx_3_422 : std_logic_vector(0 downto 0);
    signal Jr_399 : std_logic_vector(5 downto 0);
    signal R_I_424_resized : std_logic_vector(7 downto 0);
    signal R_I_424_scaled : std_logic_vector(7 downto 0);
    signal R_I_436_resized : std_logic_vector(7 downto 0);
    signal R_I_436_scaled : std_logic_vector(7 downto 0);
    signal R_I_448_resized : std_logic_vector(7 downto 0);
    signal R_I_448_scaled : std_logic_vector(7 downto 0);
    signal R_I_460_resized : std_logic_vector(7 downto 0);
    signal R_I_460_scaled : std_logic_vector(7 downto 0);
    signal R_Jr_425_resized : std_logic_vector(7 downto 0);
    signal R_Jr_425_scaled : std_logic_vector(7 downto 0);
    signal R_Jr_437_resized : std_logic_vector(7 downto 0);
    signal R_Jr_437_scaled : std_logic_vector(7 downto 0);
    signal R_Jr_449_resized : std_logic_vector(7 downto 0);
    signal R_Jr_449_scaled : std_logic_vector(7 downto 0);
    signal R_Jr_461_resized : std_logic_vector(7 downto 0);
    signal R_Jr_461_scaled : std_logic_vector(7 downto 0);
    signal ULT_u8_u1_474_wire : std_logic_vector(0 downto 0);
    signal ULT_u8_u1_480_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_426_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_426_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_426_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_438_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_450_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_word_offset_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_462_final_offset : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_index_partial_sum_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_offset_scale_factor_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_offset_scale_factor_1 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_resized_base_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_root_address : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_word_address_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_word_offset_0 : std_logic_vector(7 downto 0);
    signal aval_402 : std_logic_vector(31 downto 0);
    signal konst_376_wire_constant : std_logic_vector(7 downto 0);
    signal konst_388_wire_constant : std_logic_vector(7 downto 0);
    signal konst_405_wire_constant : std_logic_vector(1 downto 0);
    signal konst_410_wire_constant : std_logic_vector(1 downto 0);
    signal konst_415_wire_constant : std_logic_vector(1 downto 0);
    signal konst_420_wire_constant : std_logic_vector(1 downto 0);
    signal konst_473_wire_constant : std_logic_vector(7 downto 0);
    signal konst_479_wire_constant : std_logic_vector(7 downto 0);
    signal nI_378 : std_logic_vector(7 downto 0);
    signal nI_378_372_buffered : std_logic_vector(7 downto 0);
    signal nJ_390 : std_logic_vector(7 downto 0);
    signal nJ_390_384_buffered : std_logic_vector(7 downto 0);
    signal type_cast_371_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_383_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_426_offset_scale_factor_0 <= "00001000";
    array_obj_ref_426_offset_scale_factor_1 <= "00000001";
    array_obj_ref_426_resized_base_address <= "00000000";
    array_obj_ref_426_word_offset_0 <= "00000000";
    array_obj_ref_438_offset_scale_factor_0 <= "00001000";
    array_obj_ref_438_offset_scale_factor_1 <= "00000001";
    array_obj_ref_438_resized_base_address <= "00000000";
    array_obj_ref_438_word_offset_0 <= "00000000";
    array_obj_ref_450_offset_scale_factor_0 <= "00001000";
    array_obj_ref_450_offset_scale_factor_1 <= "00000001";
    array_obj_ref_450_resized_base_address <= "00000000";
    array_obj_ref_450_word_offset_0 <= "00000000";
    array_obj_ref_462_offset_scale_factor_0 <= "00001000";
    array_obj_ref_462_offset_scale_factor_1 <= "00000001";
    array_obj_ref_462_resized_base_address <= "00000000";
    array_obj_ref_462_word_offset_0 <= "00000000";
    konst_376_wire_constant <= "00000001";
    konst_388_wire_constant <= "00000001";
    konst_405_wire_constant <= "00";
    konst_410_wire_constant <= "01";
    konst_415_wire_constant <= "10";
    konst_420_wire_constant <= "11";
    konst_473_wire_constant <= "00100000";
    konst_479_wire_constant <= "00100000";
    type_cast_371_wire_constant <= "00000000";
    type_cast_383_wire_constant <= "00000000";
    phi_stmt_368: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_371_wire_constant & nI_378_372_buffered;
      req <= phi_stmt_368_req_0 & phi_stmt_368_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_368",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_368_ack_0,
          idata => idata,
          odata => I_368,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_368
    phi_stmt_380: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_383_wire_constant & nJ_390_384_buffered;
      req <= phi_stmt_380_req_0 & phi_stmt_380_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_380",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_380_ack_0,
          idata => idata,
          odata => J_380,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_380
    -- flow-through slice operator slice_394_inst
    J_idx_395 <= J_380(1 downto 0);
    slice_398_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_398_inst_req_0;
      slice_398_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_398_inst_req_1;
      slice_398_inst_ack_1<= update_ack(0);
      slice_398_inst: SliceSplitProtocol generic map(name => "slice_398_inst", in_data_width => 8, high_index => 7, low_index => 2, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => J_380, dout => Jr_399, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    nI_378_372_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_378_372_buf_req_0;
      nI_378_372_buf_ack_0<= wack(0);
      rreq(0) <= nI_378_372_buf_req_1;
      nI_378_372_buf_ack_1<= rack(0);
      nI_378_372_buf : InterlockBuffer generic map ( -- 
        name => "nI_378_372_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_378_372_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nJ_390_384_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nJ_390_384_buf_req_0;
      nJ_390_384_buf_ack_0<= wack(0);
      rreq(0) <= nJ_390_384_buf_req_1;
      nJ_390_384_buf_ack_1<= rack(0);
      nJ_390_384_buf : InterlockBuffer generic map ( -- 
        name => "nJ_390_384_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nJ_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nJ_390_384_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_426_addr_0
    process(array_obj_ref_426_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_426_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_426_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_gather_scatter
    process(aval_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := aval_402;
      ov(31 downto 0) := iv;
      array_obj_ref_426_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_index_0_resize
    process(I_368) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_368;
      ov(7 downto 0) := iv;
      R_I_424_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_index_1_rename
    process(R_Jr_425_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Jr_425_resized;
      ov(7 downto 0) := iv;
      R_Jr_425_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_index_1_resize
    process(Jr_399) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Jr_399;
      ov(5 downto 0) := iv;
      R_Jr_425_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_index_offset
    process(array_obj_ref_426_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_426_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_426_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_426_root_address_inst
    process(array_obj_ref_426_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_426_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_426_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_addr_0
    process(array_obj_ref_438_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_438_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_438_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_gather_scatter
    process(aval_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := aval_402;
      ov(31 downto 0) := iv;
      array_obj_ref_438_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_index_0_resize
    process(I_368) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_368;
      ov(7 downto 0) := iv;
      R_I_436_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_index_1_rename
    process(R_Jr_437_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Jr_437_resized;
      ov(7 downto 0) := iv;
      R_Jr_437_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_index_1_resize
    process(Jr_399) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Jr_399;
      ov(5 downto 0) := iv;
      R_Jr_437_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_index_offset
    process(array_obj_ref_438_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_438_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_438_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_438_root_address_inst
    process(array_obj_ref_438_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_438_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_438_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_addr_0
    process(array_obj_ref_450_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_450_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_450_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_gather_scatter
    process(aval_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := aval_402;
      ov(31 downto 0) := iv;
      array_obj_ref_450_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_index_0_resize
    process(I_368) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_368;
      ov(7 downto 0) := iv;
      R_I_448_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_index_1_rename
    process(R_Jr_449_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Jr_449_resized;
      ov(7 downto 0) := iv;
      R_Jr_449_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_index_1_resize
    process(Jr_399) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Jr_399;
      ov(5 downto 0) := iv;
      R_Jr_449_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_index_offset
    process(array_obj_ref_450_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_450_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_450_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_450_root_address_inst
    process(array_obj_ref_450_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_450_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_450_root_address <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_addr_0
    process(array_obj_ref_462_root_address) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_462_root_address;
      ov(7 downto 0) := iv;
      array_obj_ref_462_word_address_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_gather_scatter
    process(aval_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := aval_402;
      ov(31 downto 0) := iv;
      array_obj_ref_462_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_index_0_resize
    process(I_368) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_368;
      ov(7 downto 0) := iv;
      R_I_460_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_index_1_rename
    process(R_Jr_461_resized) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Jr_461_resized;
      ov(7 downto 0) := iv;
      R_Jr_461_scaled <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_index_1_resize
    process(Jr_399) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Jr_399;
      ov(5 downto 0) := iv;
      R_Jr_461_resized <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_index_offset
    process(array_obj_ref_462_index_partial_sum_1) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_462_index_partial_sum_1;
      ov(7 downto 0) := iv;
      array_obj_ref_462_final_offset <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_root_address_inst
    process(array_obj_ref_462_final_offset) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_462_final_offset;
      ov(7 downto 0) := iv;
      array_obj_ref_462_root_address <= ov(7 downto 0);
      --
    end process;
    if_stmt_471_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_474_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_471_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_471_branch_req_0,
          ack0 => if_stmt_471_branch_ack_0,
          ack1 => if_stmt_471_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_477_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_480_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_477_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_477_branch_req_0,
          ack0 => if_stmt_477_branch_ack_0,
          ack1 => if_stmt_477_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u8_u8_377_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= I_368;
      nI_378 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_377_inst_req_0;
      ADD_u8_u8_377_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_377_inst_req_1;
      ADD_u8_u8_377_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u8_u8_389_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= J_380;
      nJ_390 <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u8_u8_389_inst_req_0;
      ADD_u8_u8_389_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u8_u8_389_inst_req_1;
      ADD_u8_u8_389_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator EQ_u2_u1_406_inst
    process(J_idx_395) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_idx_395, konst_405_wire_constant, tmp_var);
      J_idx_0_407 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_411_inst
    process(J_idx_395) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_idx_395, konst_410_wire_constant, tmp_var);
      J_idx_1_412 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_416_inst
    process(J_idx_395) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_idx_395, konst_415_wire_constant, tmp_var);
      J_idx_2_417 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_421_inst
    process(J_idx_395) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_idx_395, konst_420_wire_constant, tmp_var);
      J_idx_3_422 <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_474_inst
    process(nJ_390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nJ_390, konst_473_wire_constant, tmp_var);
      ULT_u8_u1_474_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_480_inst
    process(nI_378) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nI_378, konst_479_wire_constant, tmp_var);
      ULT_u8_u1_480_wire <= tmp_var; --
    end process;
    -- shared split operator group (8) : array_obj_ref_426_index_0_scale array_obj_ref_438_index_0_scale array_obj_ref_450_index_0_scale array_obj_ref_462_index_0_scale 
    ApIntMul_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      data_in <= R_I_424_resized & R_I_436_resized & R_I_448_resized & R_I_460_resized;
      R_I_424_scaled <= data_out(31 downto 24);
      R_I_436_scaled <= data_out(23 downto 16);
      R_I_448_scaled <= data_out(15 downto 8);
      R_I_460_scaled <= data_out(7 downto 0);
      guard_vector(0)  <= J_idx_3_422(0);
      guard_vector(1)  <= J_idx_2_417(0);
      guard_vector(2)  <= J_idx_1_412(0);
      guard_vector(3)  <= J_idx_0_407(0);
      reqL_unguarded(3) <= array_obj_ref_426_index_0_scale_req_0;
      reqL_unguarded(2) <= array_obj_ref_438_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_450_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_462_index_0_scale_req_0;
      array_obj_ref_426_index_0_scale_ack_0 <= ackL_unguarded(3);
      array_obj_ref_438_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_450_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_462_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_426_index_0_scale_req_1;
      reqR_unguarded(2) <= array_obj_ref_438_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_450_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_462_index_0_scale_req_1;
      array_obj_ref_426_index_0_scale_ack_1 <= ackR_unguarded(3);
      array_obj_ref_438_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_450_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_462_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_8_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_8_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_8_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_8_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_8_accessRegulator_2: access_regulator_base generic map (name => "ApIntMul_group_8_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      ApIntMul_group_8_accessRegulator_3: access_regulator_base generic map (name => "ApIntMul_group_8_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      ApIntMul_group_8_gI: SplitGuardInterface generic map(name => "ApIntMul_group_8_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_8",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00001000",
          constant_width => 8,
          use_constant  => true,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 4,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_426_index_sum_1 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Jr_425_scaled & R_I_424_scaled;
      array_obj_ref_426_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <= J_idx_0_407(0);
      reqL_unguarded(0) <= array_obj_ref_426_index_sum_1_req_0;
      array_obj_ref_426_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_426_index_sum_1_req_1;
      array_obj_ref_426_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_9_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_438_index_sum_1 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Jr_437_scaled & R_I_436_scaled;
      array_obj_ref_438_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <= J_idx_1_412(0);
      reqL_unguarded(0) <= array_obj_ref_438_index_sum_1_req_0;
      array_obj_ref_438_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_438_index_sum_1_req_1;
      array_obj_ref_438_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_10_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_450_index_sum_1 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Jr_449_scaled & R_I_448_scaled;
      array_obj_ref_450_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <= J_idx_2_417(0);
      reqL_unguarded(0) <= array_obj_ref_450_index_sum_1_req_0;
      array_obj_ref_450_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_450_index_sum_1_req_1;
      array_obj_ref_450_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_462_index_sum_1 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_Jr_461_scaled & R_I_460_scaled;
      array_obj_ref_462_index_partial_sum_1 <= data_out(7 downto 0);
      guard_vector(0)  <= J_idx_3_422(0);
      reqL_unguarded(0) <= array_obj_ref_462_index_sum_1_req_0;
      array_obj_ref_462_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_462_index_sum_1_req_1;
      array_obj_ref_462_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_12_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared store operator group (0) : array_obj_ref_426_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_426_store_0_req_0;
      array_obj_ref_426_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_426_store_0_req_1;
      array_obj_ref_426_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= J_idx_0_407(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_426_word_address_0;
      data_in <= array_obj_ref_426_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(7 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : array_obj_ref_438_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_438_store_0_req_0;
      array_obj_ref_438_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_438_store_0_req_1;
      array_obj_ref_438_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= J_idx_1_412(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_438_word_address_0;
      data_in <= array_obj_ref_438_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(7 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : array_obj_ref_450_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_450_store_0_req_0;
      array_obj_ref_450_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_450_store_0_req_1;
      array_obj_ref_450_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= J_idx_2_417(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_450_word_address_0;
      data_in <= array_obj_ref_450_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(7 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : array_obj_ref_462_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(7 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_462_store_0_req_0;
      array_obj_ref_462_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_462_store_0_req_1;
      array_obj_ref_462_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= J_idx_3_422(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_462_word_address_0;
      data_in <= array_obj_ref_462_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 8,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(7 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : RPIPE_in_data_401_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_401_inst_req_0;
      RPIPE_in_data_401_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_401_inst_req_1;
      RPIPE_in_data_401_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      aval_402 <= data_out(31 downto 0);
      in_data_read_0_gI: SplitGuardInterface generic map(name => "in_data_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_read_0: InputPortRevised -- 
        generic map ( name => "in_data_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end readMatrix_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readVector is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readVector;
architecture readVector_arch of readVector is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal readVector_CP_2891_start: Boolean;
  signal readVector_CP_2891_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nI_574_493_buf_ack_1 : boolean;
  signal array_obj_ref_550_store_0_req_0 : boolean;
  signal nI_574_493_buf_req_1 : boolean;
  signal nI_574_493_buf_ack_0 : boolean;
  signal array_obj_ref_528_store_0_ack_0 : boolean;
  signal array_obj_ref_528_store_0_ack_1 : boolean;
  signal nI_574_493_buf_req_0 : boolean;
  signal array_obj_ref_528_store_0_req_0 : boolean;
  signal RPIPE_in_data_504_inst_ack_1 : boolean;
  signal RPIPE_in_data_504_inst_req_1 : boolean;
  signal array_obj_ref_528_store_0_req_1 : boolean;
  signal array_obj_ref_550_store_0_ack_0 : boolean;
  signal array_obj_ref_550_store_0_req_1 : boolean;
  signal array_obj_ref_550_store_0_ack_1 : boolean;
  signal array_obj_ref_539_store_0_ack_1 : boolean;
  signal phi_stmt_489_ack_0 : boolean;
  signal array_obj_ref_539_store_0_req_1 : boolean;
  signal phi_stmt_489_req_0 : boolean;
  signal do_while_stmt_487_branch_req_0 : boolean;
  signal phi_stmt_489_req_1 : boolean;
  signal RPIPE_in_data_504_inst_ack_0 : boolean;
  signal RPIPE_in_data_504_inst_req_0 : boolean;
  signal array_obj_ref_539_store_0_ack_0 : boolean;
  signal array_obj_ref_539_store_0_req_0 : boolean;
  signal array_obj_ref_561_store_0_req_0 : boolean;
  signal array_obj_ref_561_store_0_ack_0 : boolean;
  signal array_obj_ref_561_store_0_req_1 : boolean;
  signal array_obj_ref_561_store_0_ack_1 : boolean;
  signal do_while_stmt_487_branch_ack_0 : boolean;
  signal do_while_stmt_487_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readVector_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readVector_CP_2891_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readVector_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readVector_CP_2891_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readVector_CP_2891_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readVector_CP_2891_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readVector_CP_2891: Block -- control-path 
    signal readVector_CP_2891_elements: BooleanArray(53 downto 0);
    -- 
  begin -- 
    readVector_CP_2891_elements(0) <= readVector_CP_2891_start;
    readVector_CP_2891_symbol <= readVector_CP_2891_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_486/$entry
      -- CP-element group 0: 	 branch_block_stmt_486/do_while_stmt_487__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_486/branch_block_stmt_486__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	53 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_486/do_while_stmt_487__exit__
      -- CP-element group 1: 	 branch_block_stmt_486/$exit
      -- CP-element group 1: 	 branch_block_stmt_486/branch_block_stmt_486__exit__
      -- CP-element group 1: 	 $exit
      -- 
    readVector_CP_2891_elements(1) <= readVector_CP_2891_elements(53);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487__entry__
      -- CP-element group 2: 	 branch_block_stmt_486/do_while_stmt_487/$entry
      -- 
    readVector_CP_2891_elements(2) <= readVector_CP_2891_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	53 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487__exit__
      -- 
    -- Element group readVector_CP_2891_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_486/do_while_stmt_487/loop_back
      -- 
    -- Element group readVector_CP_2891_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	51 
    -- CP-element group 5: 	52 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_486/do_while_stmt_487/condition_done
      -- CP-element group 5: 	 branch_block_stmt_486/do_while_stmt_487/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_486/do_while_stmt_487/loop_taken/$entry
      -- 
    readVector_CP_2891_elements(5) <= readVector_CP_2891_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	50 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_486/do_while_stmt_487/loop_body_done
      -- 
    readVector_CP_2891_elements(6) <= readVector_CP_2891_elements(50);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/back_edge_to_loop_body
      -- 
    readVector_CP_2891_elements(7) <= readVector_CP_2891_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/first_time_through_loop_body
      -- 
    readVector_CP_2891_elements(8) <= readVector_CP_2891_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	49 
    -- CP-element group 9: 	29 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/$entry
      -- 
    -- Element group readVector_CP_2891_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	49 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/condition_evaluated
      -- 
    condition_evaluated_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(10), ack => do_while_stmt_487_branch_req_0); -- 
    readVector_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(15) & readVector_CP_2891_elements(49);
      gj_readVector_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/aggregated_phi_sample_req
      -- 
    readVector_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(12) & readVector_CP_2891_elements(15);
      gj_readVector_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_sample_start_
      -- 
    readVector_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(9) & readVector_CP_2891_elements(14);
      gj_readVector_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	39 
    -- CP-element group 13: 	43 
    -- CP-element group 13: 	47 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_update_start_
      -- CP-element group 13: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/aggregated_phi_update_req
      -- 
    readVector_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(9) & readVector_CP_2891_elements(35) & readVector_CP_2891_elements(39) & readVector_CP_2891_elements(43) & readVector_CP_2891_elements(47);
      gj_readVector_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	50 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_sample_completed__ps
      -- CP-element group 14: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group readVector_CP_2891_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	37 
    -- CP-element group 15: 	41 
    -- CP-element group 15: 	45 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	33 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (107) 
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_word_addrgen/root_register_ack
      -- 
    -- Element group readVector_CP_2891_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_loopback_trigger
      -- 
    readVector_CP_2891_elements(16) <= readVector_CP_2891_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_loopback_sample_req_ps
      -- CP-element group 17: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_loopback_sample_req
      -- 
    phi_stmt_489_loopback_sample_req_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_489_loopback_sample_req_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(17), ack => phi_stmt_489_req_1); -- 
    -- Element group readVector_CP_2891_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_entry_trigger
      -- 
    readVector_CP_2891_elements(18) <= readVector_CP_2891_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_entry_sample_req_ps
      -- CP-element group 19: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_entry_sample_req
      -- 
    phi_stmt_489_entry_sample_req_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_489_entry_sample_req_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(19), ack => phi_stmt_489_req_0); -- 
    -- Element group readVector_CP_2891_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_phi_mux_ack_ps
      -- CP-element group 20: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/phi_stmt_489_phi_mux_ack
      -- 
    phi_stmt_489_phi_mux_ack_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_489_ack_0, ack => readVector_CP_2891_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_sample_start__ps
      -- 
    -- Element group readVector_CP_2891_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_update_start_
      -- CP-element group 22: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_update_start__ps
      -- 
    -- Element group readVector_CP_2891_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_update_completed__ps
      -- 
    readVector_CP_2891_elements(23) <= readVector_CP_2891_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/type_cast_492_update_completed_
      -- 
    -- Element group readVector_CP_2891_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => readVector_CP_2891_elements(22), ack => readVector_CP_2891_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Sample/req
      -- CP-element group 25: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Sample/$entry
      -- 
    req_2957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(25), ack => nI_574_493_buf_req_0); -- 
    -- Element group readVector_CP_2891_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Update/req
      -- CP-element group 26: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_update_start_
      -- 
    req_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(26), ack => nI_574_493_buf_req_1); -- 
    -- Element group readVector_CP_2891_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_sample_completed_
      -- 
    ack_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_574_493_buf_ack_0, ack => readVector_CP_2891_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/R_nI_493_update_completed_
      -- 
    ack_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_574_493_buf_ack_1, ack => readVector_CP_2891_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	32 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Sample/$entry
      -- 
    rr_2972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(29), ack => RPIPE_in_data_504_inst_req_0); -- 
    readVector_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(9) & readVector_CP_2891_elements(32);
      gj_readVector_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	39 
    -- CP-element group 30: 	43 
    -- CP-element group 30: 	47 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_update_start_
      -- CP-element group 30: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Update/$entry
      -- 
    cr_2977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(30), ack => RPIPE_in_data_504_inst_req_1); -- 
    readVector_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(31) & readVector_CP_2891_elements(35) & readVector_CP_2891_elements(39) & readVector_CP_2891_elements(43) & readVector_CP_2891_elements(47);
      gj_readVector_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Sample/$exit
      -- 
    ra_2973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_504_inst_ack_0, ack => readVector_CP_2891_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32: 	41 
    -- CP-element group 32: 	45 
    -- CP-element group 32: 	33 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	29 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/RPIPE_in_data_504_update_completed_
      -- 
    ca_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_504_inst_ack_1, ack => readVector_CP_2891_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: 	32 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/array_obj_ref_528_Split/split_ack
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/array_obj_ref_528_Split/split_req
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/array_obj_ref_528_Split/$exit
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/array_obj_ref_528_Split/$entry
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/word_0/rr
      -- CP-element group 33: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/word_0/$entry
      -- 
    rr_3028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(33), ack => array_obj_ref_528_store_0_req_0); -- 
    readVector_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(15) & readVector_CP_2891_elements(32) & readVector_CP_2891_elements(35);
      gj_readVector_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/$entry
      -- CP-element group 34: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_update_start_
      -- CP-element group 34: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/word_0/cr
      -- 
    cr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(34), ack => array_obj_ref_528_store_0_req_1); -- 
    readVector_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readVector_CP_2891_elements(36);
      gj_readVector_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35: 	30 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/word_0/ra
      -- CP-element group 35: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Sample/word_access_start/word_0/$exit
      -- 
    ra_3029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_store_0_ack_0, ack => readVector_CP_2891_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	50 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_528_Update/word_access_complete/word_0/ca
      -- 
    ca_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_store_0_ack_1, ack => readVector_CP_2891_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	15 
    -- CP-element group 37: 	32 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/array_obj_ref_539_Split/$exit
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/array_obj_ref_539_Split/$entry
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/word_0/$entry
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/array_obj_ref_539_Split/split_ack
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/array_obj_ref_539_Split/split_req
      -- CP-element group 37: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/word_0/rr
      -- 
    rr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(37), ack => array_obj_ref_539_store_0_req_0); -- 
    readVector_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(15) & readVector_CP_2891_elements(32) & readVector_CP_2891_elements(39);
      gj_readVector_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_update_start_
      -- CP-element group 38: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/$entry
      -- CP-element group 38: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/word_0/$entry
      -- CP-element group 38: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/word_0/cr
      -- CP-element group 38: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/$entry
      -- 
    cr_3101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(38), ack => array_obj_ref_539_store_0_req_1); -- 
    readVector_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readVector_CP_2891_elements(40);
      gj_readVector_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	13 
    -- CP-element group 39: 	37 
    -- CP-element group 39: 	30 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/$exit
      -- CP-element group 39: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Sample/word_access_start/word_0/ra
      -- 
    ra_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_store_0_ack_0, ack => readVector_CP_2891_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	50 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/$exit
      -- CP-element group 40: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/word_access_complete/word_0/ca
      -- CP-element group 40: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_539_Update/$exit
      -- 
    ca_3102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_store_0_ack_1, ack => readVector_CP_2891_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	15 
    -- CP-element group 41: 	32 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/array_obj_ref_550_Split/split_ack
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/array_obj_ref_550_Split/split_req
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/array_obj_ref_550_Split/$entry
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/array_obj_ref_550_Split/$exit
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/$entry
      -- 
    rr_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(41), ack => array_obj_ref_550_store_0_req_0); -- 
    readVector_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(15) & readVector_CP_2891_elements(32) & readVector_CP_2891_elements(43);
      gj_readVector_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/word_0/cr
      -- CP-element group 42: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/$entry
      -- CP-element group 42: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_update_start_
      -- 
    cr_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(42), ack => array_obj_ref_550_store_0_req_1); -- 
    readVector_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readVector_CP_2891_elements(44);
      gj_readVector_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	13 
    -- CP-element group 43: 	41 
    -- CP-element group 43: 	30 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/word_0/ra
      -- CP-element group 43: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Sample/$exit
      -- 
    ra_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_550_store_0_ack_0, ack => readVector_CP_2891_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_550_update_completed_
      -- 
    ca_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_550_store_0_ack_1, ack => readVector_CP_2891_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	15 
    -- CP-element group 45: 	32 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/array_obj_ref_561_Split/$entry
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/array_obj_ref_561_Split/$exit
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/array_obj_ref_561_Split/split_req
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/array_obj_ref_561_Split/split_ack
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/$entry
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/word_0/rr
      -- 
    rr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(45), ack => array_obj_ref_561_store_0_req_0); -- 
    readVector_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(15) & readVector_CP_2891_elements(32) & readVector_CP_2891_elements(47);
      gj_readVector_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_update_start_
      -- CP-element group 46: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/$entry
      -- CP-element group 46: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/word_0/cr
      -- 
    cr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readVector_CP_2891_elements(46), ack => array_obj_ref_561_store_0_req_1); -- 
    readVector_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readVector_CP_2891_elements(48);
      gj_readVector_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	13 
    -- CP-element group 47: 	45 
    -- CP-element group 47: 	30 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Sample/word_access_start/word_0/ra
      -- 
    ra_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_store_0_ack_0, ack => readVector_CP_2891_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/array_obj_ref_561_Update/word_access_complete/word_0/ca
      -- 
    ca_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_store_0_ack_1, ack => readVector_CP_2891_elements(48)); -- 
    -- CP-element group 49:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	9 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	10 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group readVector_CP_2891_elements(49) is a control-delay.
    cp_element_49_delay: control_delay_element  generic map(name => " 49_delay", delay_value => 1)  port map(req => readVector_CP_2891_elements(9), ack => readVector_CP_2891_elements(49), clk => clk, reset =>reset);
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	14 
    -- CP-element group 50: 	36 
    -- CP-element group 50: 	40 
    -- CP-element group 50: 	44 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	6 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_486/do_while_stmt_487/do_while_stmt_487_loop_body/$exit
      -- 
    readVector_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "readVector_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= readVector_CP_2891_elements(14) & readVector_CP_2891_elements(36) & readVector_CP_2891_elements(40) & readVector_CP_2891_elements(44) & readVector_CP_2891_elements(48);
      gj_readVector_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readVector_CP_2891_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	5 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_486/do_while_stmt_487/loop_exit/$exit
      -- CP-element group 51: 	 branch_block_stmt_486/do_while_stmt_487/loop_exit/ack
      -- 
    ack_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_487_branch_ack_0, ack => readVector_CP_2891_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	5 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_486/do_while_stmt_487/loop_taken/$exit
      -- CP-element group 52: 	 branch_block_stmt_486/do_while_stmt_487/loop_taken/ack
      -- 
    ack_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_487_branch_ack_1, ack => readVector_CP_2891_elements(52)); -- 
    -- CP-element group 53:  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	3 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	1 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_486/do_while_stmt_487/$exit
      -- 
    readVector_CP_2891_elements(53) <= readVector_CP_2891_elements(3);
    readVector_do_while_stmt_487_terminator_3236: loop_terminator -- 
      generic map (name => " readVector_do_while_stmt_487_terminator_3236", max_iterations_in_flight =>7) 
      port map(loop_body_exit => readVector_CP_2891_elements(6),loop_continue => readVector_CP_2891_elements(52),loop_terminate => readVector_CP_2891_elements(51),loop_back => readVector_CP_2891_elements(4),loop_exit => readVector_CP_2891_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_489_phi_seq_2964_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= readVector_CP_2891_elements(18);
      readVector_CP_2891_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= readVector_CP_2891_elements(21);
      readVector_CP_2891_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= readVector_CP_2891_elements(23);
      readVector_CP_2891_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= readVector_CP_2891_elements(16);
      readVector_CP_2891_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= readVector_CP_2891_elements(27);
      readVector_CP_2891_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= readVector_CP_2891_elements(28);
      readVector_CP_2891_elements(17) <= phi_mux_reqs(1);
      phi_stmt_489_phi_seq_2964 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_489_phi_seq_2964") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => readVector_CP_2891_elements(11), 
          phi_sample_ack => readVector_CP_2891_elements(14), 
          phi_update_req => readVector_CP_2891_elements(13), 
          phi_update_ack => readVector_CP_2891_elements(15), 
          phi_mux_ack => readVector_CP_2891_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2916_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= readVector_CP_2891_elements(7);
        preds(1)  <= readVector_CP_2891_elements(8);
        entry_tmerge_2916 : transition_merge -- 
          generic map(name => " entry_tmerge_2916")
          port map (preds => preds, symbol_out => readVector_CP_2891_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_489 : std_logic_vector(7 downto 0);
    signal I_idx_0_510 : std_logic_vector(0 downto 0);
    signal I_idx_1_515 : std_logic_vector(0 downto 0);
    signal I_idx_2_520 : std_logic_vector(0 downto 0);
    signal I_idx_3_525 : std_logic_vector(0 downto 0);
    signal I_idx_498 : std_logic_vector(1 downto 0);
    signal Ir_502 : std_logic_vector(5 downto 0);
    signal R_Ir_527_resized : std_logic_vector(2 downto 0);
    signal R_Ir_527_scaled : std_logic_vector(2 downto 0);
    signal R_Ir_538_resized : std_logic_vector(2 downto 0);
    signal R_Ir_538_scaled : std_logic_vector(2 downto 0);
    signal R_Ir_549_resized : std_logic_vector(2 downto 0);
    signal R_Ir_549_scaled : std_logic_vector(2 downto 0);
    signal R_Ir_560_resized : std_logic_vector(2 downto 0);
    signal R_Ir_560_scaled : std_logic_vector(2 downto 0);
    signal ULT_u8_u1_578_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_528_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_528_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_528_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_528_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_528_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_528_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_528_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_539_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_539_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_550_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_550_word_offset_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_561_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_561_word_offset_0 : std_logic_vector(2 downto 0);
    signal konst_508_wire_constant : std_logic_vector(1 downto 0);
    signal konst_513_wire_constant : std_logic_vector(1 downto 0);
    signal konst_518_wire_constant : std_logic_vector(1 downto 0);
    signal konst_523_wire_constant : std_logic_vector(1 downto 0);
    signal konst_572_wire_constant : std_logic_vector(7 downto 0);
    signal konst_577_wire_constant : std_logic_vector(7 downto 0);
    signal nI_574 : std_logic_vector(7 downto 0);
    signal nI_574_493_buffered : std_logic_vector(7 downto 0);
    signal temp_val_505 : std_logic_vector(31 downto 0);
    signal type_cast_492_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_528_offset_scale_factor_0 <= "001";
    array_obj_ref_528_resized_base_address <= "000";
    array_obj_ref_528_word_offset_0 <= "000";
    array_obj_ref_539_offset_scale_factor_0 <= "001";
    array_obj_ref_539_resized_base_address <= "000";
    array_obj_ref_539_word_offset_0 <= "000";
    array_obj_ref_550_offset_scale_factor_0 <= "001";
    array_obj_ref_550_resized_base_address <= "000";
    array_obj_ref_550_word_offset_0 <= "000";
    array_obj_ref_561_offset_scale_factor_0 <= "001";
    array_obj_ref_561_resized_base_address <= "000";
    array_obj_ref_561_word_offset_0 <= "000";
    konst_508_wire_constant <= "00";
    konst_513_wire_constant <= "01";
    konst_518_wire_constant <= "10";
    konst_523_wire_constant <= "11";
    konst_572_wire_constant <= "00000001";
    konst_577_wire_constant <= "00100000";
    type_cast_492_wire_constant <= "00000000";
    phi_stmt_489: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_492_wire_constant & nI_574_493_buffered;
      req <= phi_stmt_489_req_0 & phi_stmt_489_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_489",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_489_ack_0,
          idata => idata,
          odata => I_489,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_489
    -- flow-through slice operator slice_497_inst
    I_idx_498 <= I_489(1 downto 0);
    -- flow-through slice operator slice_501_inst
    Ir_502 <= I_489(7 downto 2);
    nI_574_493_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_574_493_buf_req_0;
      nI_574_493_buf_ack_0<= wack(0);
      rreq(0) <= nI_574_493_buf_req_1;
      nI_574_493_buf_ack_1<= rack(0);
      nI_574_493_buf : InterlockBuffer generic map ( -- 
        name => "nI_574_493_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_574_493_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_528_addr_0
    process(array_obj_ref_528_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_528_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_528_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_528_gather_scatter
    process(temp_val_505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := temp_val_505;
      ov(31 downto 0) := iv;
      array_obj_ref_528_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_528_index_0_rename
    process(R_Ir_527_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_527_resized;
      ov(2 downto 0) := iv;
      R_Ir_527_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_528_index_0_resize
    process(Ir_502) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Ir_502;
      ov := iv(2 downto 0);
      R_Ir_527_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_528_index_offset
    process(R_Ir_527_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_527_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_528_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_528_root_address_inst
    process(array_obj_ref_528_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_528_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_528_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_addr_0
    process(array_obj_ref_539_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_539_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_539_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_gather_scatter
    process(temp_val_505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := temp_val_505;
      ov(31 downto 0) := iv;
      array_obj_ref_539_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_index_0_rename
    process(R_Ir_538_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_538_resized;
      ov(2 downto 0) := iv;
      R_Ir_538_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_index_0_resize
    process(Ir_502) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Ir_502;
      ov := iv(2 downto 0);
      R_Ir_538_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_index_offset
    process(R_Ir_538_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_538_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_539_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_539_root_address_inst
    process(array_obj_ref_539_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_539_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_539_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_addr_0
    process(array_obj_ref_550_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_550_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_550_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_gather_scatter
    process(temp_val_505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := temp_val_505;
      ov(31 downto 0) := iv;
      array_obj_ref_550_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_index_0_rename
    process(R_Ir_549_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_549_resized;
      ov(2 downto 0) := iv;
      R_Ir_549_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_index_0_resize
    process(Ir_502) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Ir_502;
      ov := iv(2 downto 0);
      R_Ir_549_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_index_offset
    process(R_Ir_549_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_549_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_550_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_550_root_address_inst
    process(array_obj_ref_550_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_550_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_550_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_addr_0
    process(array_obj_ref_561_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_561_root_address;
      ov(2 downto 0) := iv;
      array_obj_ref_561_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_gather_scatter
    process(temp_val_505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := temp_val_505;
      ov(31 downto 0) := iv;
      array_obj_ref_561_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_index_0_rename
    process(R_Ir_560_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_560_resized;
      ov(2 downto 0) := iv;
      R_Ir_560_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_index_0_resize
    process(Ir_502) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := Ir_502;
      ov := iv(2 downto 0);
      R_Ir_560_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_index_offset
    process(R_Ir_560_scaled) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_Ir_560_scaled;
      ov(2 downto 0) := iv;
      array_obj_ref_561_final_offset <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_561_root_address_inst
    process(array_obj_ref_561_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_561_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_561_root_address <= ov(2 downto 0);
      --
    end process;
    do_while_stmt_487_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_578_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_487_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_487_branch_req_0,
          ack0 => do_while_stmt_487_branch_ack_0,
          ack1 => do_while_stmt_487_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u8_u8_573_inst
    process(I_489) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_489, konst_572_wire_constant, tmp_var);
      nI_574 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_509_inst
    process(I_idx_498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_idx_498, konst_508_wire_constant, tmp_var);
      I_idx_0_510 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_514_inst
    process(I_idx_498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_idx_498, konst_513_wire_constant, tmp_var);
      I_idx_1_515 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_519_inst
    process(I_idx_498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_idx_498, konst_518_wire_constant, tmp_var);
      I_idx_2_520 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_524_inst
    process(I_idx_498) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_idx_498, konst_523_wire_constant, tmp_var);
      I_idx_3_525 <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_578_inst
    process(nI_574) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nI_574, konst_577_wire_constant, tmp_var);
      ULT_u8_u1_578_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_528_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_528_store_0_req_0;
      array_obj_ref_528_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_528_store_0_req_1;
      array_obj_ref_528_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= I_idx_0_510(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_528_word_address_0;
      data_in <= array_obj_ref_528_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(2 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : array_obj_ref_539_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_539_store_0_req_0;
      array_obj_ref_539_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_539_store_0_req_1;
      array_obj_ref_539_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= I_idx_1_515(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_539_word_address_0;
      data_in <= array_obj_ref_539_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(2 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : array_obj_ref_550_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_550_store_0_req_0;
      array_obj_ref_550_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_550_store_0_req_1;
      array_obj_ref_550_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= I_idx_2_520(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_550_word_address_0;
      data_in <= array_obj_ref_550_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(2 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : array_obj_ref_561_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_561_store_0_req_0;
      array_obj_ref_561_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_561_store_0_req_1;
      array_obj_ref_561_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= I_idx_3_525(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_561_word_address_0;
      data_in <= array_obj_ref_561_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(2 downto 0),
          mdata => memory_space_7_sr_data(31 downto 0),
          mtag => memory_space_7_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : RPIPE_in_data_504_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_504_inst_req_0;
      RPIPE_in_data_504_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_504_inst_req_1;
      RPIPE_in_data_504_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      temp_val_505 <= data_out(31 downto 0);
      in_data_read_0_gI: SplitGuardInterface generic map(name => "in_data_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_read_0: InputPortRevised -- 
        generic map ( name => "in_data_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end readVector_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendVector is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(4 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendVector;
architecture sendVector_arch of sendVector is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendVector_CP_3237_start: Boolean;
  signal sendVector_CP_3237_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nI_599_589_buf_ack_1 : boolean;
  signal nI_599_589_buf_req_1 : boolean;
  signal WPIPE_out_data_591_inst_req_1 : boolean;
  signal WPIPE_out_data_591_inst_ack_1 : boolean;
  signal do_while_stmt_583_branch_ack_0 : boolean;
  signal WPIPE_out_data_591_inst_req_0 : boolean;
  signal WPIPE_out_data_591_inst_ack_0 : boolean;
  signal array_obj_ref_593_load_0_req_0 : boolean;
  signal nI_599_589_buf_req_0 : boolean;
  signal do_while_stmt_583_branch_ack_1 : boolean;
  signal nI_599_589_buf_ack_0 : boolean;
  signal array_obj_ref_593_load_0_ack_0 : boolean;
  signal array_obj_ref_593_load_0_ack_1 : boolean;
  signal array_obj_ref_593_load_0_req_1 : boolean;
  signal do_while_stmt_583_branch_req_0 : boolean;
  signal phi_stmt_585_req_1 : boolean;
  signal phi_stmt_585_req_0 : boolean;
  signal phi_stmt_585_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendVector_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendVector_CP_3237_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendVector_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendVector_CP_3237_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendVector_CP_3237_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendVector_CP_3237_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendVector_CP_3237: Block -- control-path 
    signal sendVector_CP_3237_elements: BooleanArray(40 downto 0);
    -- 
  begin -- 
    sendVector_CP_3237_elements(0) <= sendVector_CP_3237_start;
    sendVector_CP_3237_symbol <= sendVector_CP_3237_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_582/$entry
      -- CP-element group 0: 	 branch_block_stmt_582/branch_block_stmt_582__entry__
      -- CP-element group 0: 	 branch_block_stmt_582/do_while_stmt_583__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	40 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_582/$exit
      -- CP-element group 1: 	 branch_block_stmt_582/branch_block_stmt_582__exit__
      -- CP-element group 1: 	 branch_block_stmt_582/do_while_stmt_583__exit__
      -- 
    sendVector_CP_3237_elements(1) <= sendVector_CP_3237_elements(40);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_582/do_while_stmt_583/$entry
      -- CP-element group 2: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583__entry__
      -- 
    sendVector_CP_3237_elements(2) <= sendVector_CP_3237_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	40 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583__exit__
      -- 
    -- Element group sendVector_CP_3237_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_582/do_while_stmt_583/loop_back
      -- 
    -- Element group sendVector_CP_3237_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	38 
    -- CP-element group 5: 	39 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_582/do_while_stmt_583/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_582/do_while_stmt_583/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_582/do_while_stmt_583/condition_done
      -- 
    sendVector_CP_3237_elements(5) <= sendVector_CP_3237_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	37 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_582/do_while_stmt_583/loop_body_done
      -- 
    sendVector_CP_3237_elements(6) <= sendVector_CP_3237_elements(37);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/back_edge_to_loop_body
      -- 
    sendVector_CP_3237_elements(7) <= sendVector_CP_3237_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/first_time_through_loop_body
      -- 
    sendVector_CP_3237_elements(8) <= sendVector_CP_3237_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	36 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/loop_body_start
      -- 
    -- Element group sendVector_CP_3237_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	36 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/condition_evaluated
      -- 
    condition_evaluated_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(10), ack => do_while_stmt_583_branch_req_0); -- 
    sendVector_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(15) & sendVector_CP_3237_elements(36);
      gj_sendVector_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_sample_start__ps
      -- 
    sendVector_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(12) & sendVector_CP_3237_elements(15);
      gj_sendVector_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_sample_start_
      -- 
    sendVector_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(9) & sendVector_CP_3237_elements(14);
      gj_sendVector_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	31 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_update_start_
      -- CP-element group 13: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_update_start__ps
      -- 
    sendVector_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(9) & sendVector_CP_3237_elements(31);
      gj_sendVector_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_sample_completed__ps
      -- 
    -- Element group sendVector_CP_3237_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	29 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (29) 
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_final_index_sum_regn/req
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_update_completed__ps
      -- 
    -- Element group sendVector_CP_3237_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_loopback_trigger
      -- 
    sendVector_CP_3237_elements(16) <= sendVector_CP_3237_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_loopback_sample_req_ps
      -- 
    phi_stmt_585_loopback_sample_req_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_loopback_sample_req_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(17), ack => phi_stmt_585_req_1); -- 
    -- Element group sendVector_CP_3237_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_entry_trigger
      -- 
    sendVector_CP_3237_elements(18) <= sendVector_CP_3237_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_entry_sample_req_ps
      -- 
    phi_stmt_585_entry_sample_req_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_entry_sample_req_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(19), ack => phi_stmt_585_req_0); -- 
    -- Element group sendVector_CP_3237_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/phi_stmt_585_phi_mux_ack_ps
      -- 
    phi_stmt_585_phi_mux_ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_585_ack_0, ack => sendVector_CP_3237_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_sample_completed_
      -- 
    -- Element group sendVector_CP_3237_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_update_start_
      -- 
    -- Element group sendVector_CP_3237_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_update_completed__ps
      -- 
    sendVector_CP_3237_elements(23) <= sendVector_CP_3237_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/type_cast_588_update_completed_
      -- 
    -- Element group sendVector_CP_3237_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => sendVector_CP_3237_elements(22), ack => sendVector_CP_3237_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Sample/req
      -- CP-element group 25: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_sample_start_
      -- 
    req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(25), ack => nI_599_589_buf_req_0); -- 
    -- Element group sendVector_CP_3237_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Update/req
      -- CP-element group 26: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_update_start_
      -- 
    req_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(26), ack => nI_599_589_buf_req_1); -- 
    -- Element group sendVector_CP_3237_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_sample_completed_
      -- 
    ack_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_599_589_buf_ack_0, ack => sendVector_CP_3237_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/R_nI_589_update_completed_
      -- 
    ack_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_599_589_buf_ack_1, ack => sendVector_CP_3237_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/word_0/rr
      -- CP-element group 29: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/$entry
      -- 
    rr_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(29), ack => array_obj_ref_593_load_0_req_0); -- 
    sendVector_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(15) & sendVector_CP_3237_elements(31);
      gj_sendVector_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	34 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/word_0/$entry
      -- CP-element group 30: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_update_start_
      -- CP-element group 30: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/$entry
      -- CP-element group 30: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/word_0/cr
      -- CP-element group 30: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/$entry
      -- 
    cr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(30), ack => array_obj_ref_593_load_0_req_1); -- 
    sendVector_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendVector_CP_3237_elements(34);
      gj_sendVector_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Sample/word_access_start/word_0/ra
      -- 
    ra_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_593_load_0_ack_0, ack => sendVector_CP_3237_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/array_obj_ref_593_Merge/merge_ack
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/array_obj_ref_593_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/array_obj_ref_593_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/array_obj_ref_593_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/array_obj_ref_593_Update/$exit
      -- 
    ca_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_593_load_0_ack_1, ack => sendVector_CP_3237_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_sample_start_
      -- 
    req_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(33), ack => WPIPE_out_data_591_inst_req_0); -- 
    sendVector_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(32) & sendVector_CP_3237_elements(35);
      gj_sendVector_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	30 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Update/req
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_update_start_
      -- CP-element group 34: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_sample_completed_
      -- 
    ack_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_591_inst_ack_0, ack => sendVector_CP_3237_elements(34)); -- 
    req_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendVector_CP_3237_elements(34), ack => WPIPE_out_data_591_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/WPIPE_out_data_591_update_completed_
      -- 
    ack_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_591_inst_ack_1, ack => sendVector_CP_3237_elements(35)); -- 
    -- CP-element group 36:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	10 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendVector_CP_3237_elements(36) is a control-delay.
    cp_element_36_delay: control_delay_element  generic map(name => " 36_delay", delay_value => 1)  port map(req => sendVector_CP_3237_elements(9), ack => sendVector_CP_3237_elements(36), clk => clk, reset =>reset);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	6 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_582/do_while_stmt_583/do_while_stmt_583_loop_body/$exit
      -- 
    sendVector_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendVector_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendVector_CP_3237_elements(14) & sendVector_CP_3237_elements(35);
      gj_sendVector_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendVector_CP_3237_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_582/do_while_stmt_583/loop_exit/$exit
      -- CP-element group 38: 	 branch_block_stmt_582/do_while_stmt_583/loop_exit/ack
      -- 
    ack_3392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_583_branch_ack_0, ack => sendVector_CP_3237_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	5 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_582/do_while_stmt_583/loop_taken/$exit
      -- CP-element group 39: 	 branch_block_stmt_582/do_while_stmt_583/loop_taken/ack
      -- 
    ack_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_583_branch_ack_1, ack => sendVector_CP_3237_elements(39)); -- 
    -- CP-element group 40:  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	3 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	1 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_582/do_while_stmt_583/$exit
      -- 
    sendVector_CP_3237_elements(40) <= sendVector_CP_3237_elements(3);
    sendVector_do_while_stmt_583_terminator_3397: loop_terminator -- 
      generic map (name => " sendVector_do_while_stmt_583_terminator_3397", max_iterations_in_flight =>7) 
      port map(loop_body_exit => sendVector_CP_3237_elements(6),loop_continue => sendVector_CP_3237_elements(39),loop_terminate => sendVector_CP_3237_elements(38),loop_back => sendVector_CP_3237_elements(4),loop_exit => sendVector_CP_3237_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_585_phi_seq_3310_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendVector_CP_3237_elements(18);
      sendVector_CP_3237_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendVector_CP_3237_elements(21);
      sendVector_CP_3237_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= sendVector_CP_3237_elements(23);
      sendVector_CP_3237_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= sendVector_CP_3237_elements(16);
      sendVector_CP_3237_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendVector_CP_3237_elements(27);
      sendVector_CP_3237_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= sendVector_CP_3237_elements(28);
      sendVector_CP_3237_elements(17) <= phi_mux_reqs(1);
      phi_stmt_585_phi_seq_3310 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_585_phi_seq_3310") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendVector_CP_3237_elements(11), 
          phi_sample_ack => sendVector_CP_3237_elements(14), 
          phi_update_req => sendVector_CP_3237_elements(13), 
          phi_update_ack => sendVector_CP_3237_elements(15), 
          phi_mux_ack => sendVector_CP_3237_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3262_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendVector_CP_3237_elements(7);
        preds(1)  <= sendVector_CP_3237_elements(8);
        entry_tmerge_3262 : transition_merge -- 
          generic map(name => " entry_tmerge_3262")
          port map (preds => preds, symbol_out => sendVector_CP_3237_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_585 : std_logic_vector(7 downto 0);
    signal R_I_592_resized : std_logic_vector(4 downto 0);
    signal R_I_592_scaled : std_logic_vector(4 downto 0);
    signal ULT_u8_u1_603_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_593_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_593_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_593_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_593_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_593_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_593_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_593_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_593_word_offset_0 : std_logic_vector(4 downto 0);
    signal konst_597_wire_constant : std_logic_vector(7 downto 0);
    signal konst_602_wire_constant : std_logic_vector(7 downto 0);
    signal nI_599 : std_logic_vector(7 downto 0);
    signal nI_599_589_buffered : std_logic_vector(7 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_593_offset_scale_factor_0 <= "00001";
    array_obj_ref_593_resized_base_address <= "00000";
    array_obj_ref_593_word_offset_0 <= "00000";
    konst_597_wire_constant <= "00000001";
    konst_602_wire_constant <= "00100000";
    type_cast_588_wire_constant <= "00000000";
    phi_stmt_585: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_588_wire_constant & nI_599_589_buffered;
      req <= phi_stmt_585_req_0 & phi_stmt_585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_585",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_585_ack_0,
          idata => idata,
          odata => I_585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_585
    nI_599_589_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_599_589_buf_req_0;
      nI_599_589_buf_ack_0<= wack(0);
      rreq(0) <= nI_599_589_buf_req_1;
      nI_599_589_buf_ack_1<= rack(0);
      nI_599_589_buf : InterlockBuffer generic map ( -- 
        name => "nI_599_589_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_599_589_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_593_addr_0
    process(array_obj_ref_593_root_address) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_593_root_address;
      ov(4 downto 0) := iv;
      array_obj_ref_593_word_address_0 <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_gather_scatter
    process(array_obj_ref_593_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_593_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_593_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_index_0_rename
    process(R_I_592_resized) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_592_resized;
      ov(4 downto 0) := iv;
      R_I_592_scaled <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_index_0_resize
    process(I_585) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_585;
      ov := iv(4 downto 0);
      R_I_592_resized <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_index_offset
    process(R_I_592_scaled) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_592_scaled;
      ov(4 downto 0) := iv;
      array_obj_ref_593_final_offset <= ov(4 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_593_root_address_inst
    process(array_obj_ref_593_final_offset) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(4 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_593_final_offset;
      ov(4 downto 0) := iv;
      array_obj_ref_593_root_address <= ov(4 downto 0);
      --
    end process;
    do_while_stmt_583_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u8_u1_603_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_583_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_583_branch_req_0,
          ack0 => do_while_stmt_583_branch_ack_0,
          ack1 => do_while_stmt_583_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u8_u8_598_inst
    process(I_585) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_585, konst_597_wire_constant, tmp_var);
      nI_599 <= tmp_var; --
    end process;
    -- binary operator ULT_u8_u1_603_inst
    process(nI_599) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(nI_599, konst_602_wire_constant, tmp_var);
      ULT_u8_u1_603_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_593_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_593_load_0_req_0;
      array_obj_ref_593_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_593_load_0_req_1;
      array_obj_ref_593_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_593_word_address_0;
      array_obj_ref_593_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 5,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(4 downto 0),
          mtag => memory_space_8_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(31 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_out_data_591_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_591_inst_req_0;
      WPIPE_out_data_591_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_591_inst_req_1;
      WPIPE_out_data_591_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= array_obj_ref_593_wire;
      out_data_write_0_gI: SplitGuardInterface generic map(name => "out_data_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_write_0: OutputPortRevised -- 
        generic map ( name => "out_data", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendVector_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(15 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(15 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(15 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(15 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(5 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(5 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(5 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(5 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(35 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(4 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module dotP_even
  component dotP_even is -- 
    generic (tag_length : integer); 
    port ( -- 
      R : in  std_logic_vector(7 downto 0);
      result : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module dotP_even
  signal dotP_even_R :  std_logic_vector(7 downto 0);
  signal dotP_even_result :  std_logic_vector(31 downto 0);
  signal dotP_even_in_args    : std_logic_vector(7 downto 0);
  signal dotP_even_out_args   : std_logic_vector(31 downto 0);
  signal dotP_even_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal dotP_even_tag_out   : std_logic_vector(1 downto 0);
  signal dotP_even_start_req : std_logic;
  signal dotP_even_start_ack : std_logic;
  signal dotP_even_fin_req   : std_logic;
  signal dotP_even_fin_ack : std_logic;
  -- caller side aggregated signals for module dotP_even
  signal dotP_even_call_reqs: std_logic_vector(0 downto 0);
  signal dotP_even_call_acks: std_logic_vector(0 downto 0);
  signal dotP_even_return_reqs: std_logic_vector(0 downto 0);
  signal dotP_even_return_acks: std_logic_vector(0 downto 0);
  signal dotP_even_call_data: std_logic_vector(7 downto 0);
  signal dotP_even_call_tag: std_logic_vector(0 downto 0);
  signal dotP_even_return_data: std_logic_vector(31 downto 0);
  signal dotP_even_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module dotP_odd
  component dotP_odd is -- 
    generic (tag_length : integer); 
    port ( -- 
      R : in  std_logic_vector(7 downto 0);
      result : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module dotP_odd
  signal dotP_odd_R :  std_logic_vector(7 downto 0);
  signal dotP_odd_result :  std_logic_vector(31 downto 0);
  signal dotP_odd_in_args    : std_logic_vector(7 downto 0);
  signal dotP_odd_out_args   : std_logic_vector(31 downto 0);
  signal dotP_odd_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal dotP_odd_tag_out   : std_logic_vector(1 downto 0);
  signal dotP_odd_start_req : std_logic;
  signal dotP_odd_start_ack : std_logic;
  signal dotP_odd_fin_req   : std_logic;
  signal dotP_odd_fin_ack : std_logic;
  -- caller side aggregated signals for module dotP_odd
  signal dotP_odd_call_reqs: std_logic_vector(0 downto 0);
  signal dotP_odd_call_acks: std_logic_vector(0 downto 0);
  signal dotP_odd_return_reqs: std_logic_vector(0 downto 0);
  signal dotP_odd_return_acks: std_logic_vector(0 downto 0);
  signal dotP_odd_call_data: std_logic_vector(7 downto 0);
  signal dotP_odd_call_tag: std_logic_vector(0 downto 0);
  signal dotP_odd_return_data: std_logic_vector(31 downto 0);
  signal dotP_odd_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module multiplyMatrixVector
  component multiplyMatrixVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      dotP_even_call_reqs : out  std_logic_vector(0 downto 0);
      dotP_even_call_acks : in   std_logic_vector(0 downto 0);
      dotP_even_call_data : out  std_logic_vector(7 downto 0);
      dotP_even_call_tag  :  out  std_logic_vector(0 downto 0);
      dotP_even_return_reqs : out  std_logic_vector(0 downto 0);
      dotP_even_return_acks : in   std_logic_vector(0 downto 0);
      dotP_even_return_data : in   std_logic_vector(31 downto 0);
      dotP_even_return_tag :  in   std_logic_vector(0 downto 0);
      dotP_odd_call_reqs : out  std_logic_vector(0 downto 0);
      dotP_odd_call_acks : in   std_logic_vector(0 downto 0);
      dotP_odd_call_data : out  std_logic_vector(7 downto 0);
      dotP_odd_call_tag  :  out  std_logic_vector(0 downto 0);
      dotP_odd_return_reqs : out  std_logic_vector(0 downto 0);
      dotP_odd_return_acks : in   std_logic_vector(0 downto 0);
      dotP_odd_return_data : in   std_logic_vector(31 downto 0);
      dotP_odd_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module multiplyMatrixVector
  signal multiplyMatrixVector_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal multiplyMatrixVector_tag_out   : std_logic_vector(1 downto 0);
  signal multiplyMatrixVector_start_req : std_logic;
  signal multiplyMatrixVector_start_ack : std_logic;
  signal multiplyMatrixVector_fin_req   : std_logic;
  signal multiplyMatrixVector_fin_ack : std_logic;
  -- caller side aggregated signals for module multiplyMatrixVector
  signal multiplyMatrixVector_call_reqs: std_logic_vector(0 downto 0);
  signal multiplyMatrixVector_call_acks: std_logic_vector(0 downto 0);
  signal multiplyMatrixVector_return_reqs: std_logic_vector(0 downto 0);
  signal multiplyMatrixVector_return_acks: std_logic_vector(0 downto 0);
  signal multiplyMatrixVector_call_tag: std_logic_vector(0 downto 0);
  signal multiplyMatrixVector_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module mvp_daemon
  component mvp_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      readVector_call_reqs : out  std_logic_vector(0 downto 0);
      readVector_call_acks : in   std_logic_vector(0 downto 0);
      readVector_call_tag  :  out  std_logic_vector(0 downto 0);
      readVector_return_reqs : out  std_logic_vector(0 downto 0);
      readVector_return_acks : in   std_logic_vector(0 downto 0);
      readVector_return_tag :  in   std_logic_vector(0 downto 0);
      multiplyMatrixVector_call_reqs : out  std_logic_vector(0 downto 0);
      multiplyMatrixVector_call_acks : in   std_logic_vector(0 downto 0);
      multiplyMatrixVector_call_tag  :  out  std_logic_vector(0 downto 0);
      multiplyMatrixVector_return_reqs : out  std_logic_vector(0 downto 0);
      multiplyMatrixVector_return_acks : in   std_logic_vector(0 downto 0);
      multiplyMatrixVector_return_tag :  in   std_logic_vector(0 downto 0);
      readMatrix_call_reqs : out  std_logic_vector(0 downto 0);
      readMatrix_call_acks : in   std_logic_vector(0 downto 0);
      readMatrix_call_tag  :  out  std_logic_vector(0 downto 0);
      readMatrix_return_reqs : out  std_logic_vector(0 downto 0);
      readMatrix_return_acks : in   std_logic_vector(0 downto 0);
      readMatrix_return_tag :  in   std_logic_vector(0 downto 0);
      sendVector_call_reqs : out  std_logic_vector(0 downto 0);
      sendVector_call_acks : in   std_logic_vector(0 downto 0);
      sendVector_call_tag  :  out  std_logic_vector(0 downto 0);
      sendVector_return_reqs : out  std_logic_vector(0 downto 0);
      sendVector_return_acks : in   std_logic_vector(0 downto 0);
      sendVector_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module mvp_daemon
  signal mvp_daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal mvp_daemon_tag_out   : std_logic_vector(1 downto 0);
  signal mvp_daemon_start_req : std_logic;
  signal mvp_daemon_start_ack : std_logic;
  signal mvp_daemon_fin_req   : std_logic;
  signal mvp_daemon_fin_ack : std_logic;
  -- declarations related to module readMatrix
  component readMatrix is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readMatrix
  signal readMatrix_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readMatrix_tag_out   : std_logic_vector(1 downto 0);
  signal readMatrix_start_req : std_logic;
  signal readMatrix_start_ack : std_logic;
  signal readMatrix_fin_req   : std_logic;
  signal readMatrix_fin_ack : std_logic;
  -- caller side aggregated signals for module readMatrix
  signal readMatrix_call_reqs: std_logic_vector(0 downto 0);
  signal readMatrix_call_acks: std_logic_vector(0 downto 0);
  signal readMatrix_return_reqs: std_logic_vector(0 downto 0);
  signal readMatrix_return_acks: std_logic_vector(0 downto 0);
  signal readMatrix_call_tag: std_logic_vector(0 downto 0);
  signal readMatrix_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module readVector
  component readVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readVector
  signal readVector_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readVector_tag_out   : std_logic_vector(1 downto 0);
  signal readVector_start_req : std_logic;
  signal readVector_start_ack : std_logic;
  signal readVector_fin_req   : std_logic;
  signal readVector_fin_ack : std_logic;
  -- caller side aggregated signals for module readVector
  signal readVector_call_reqs: std_logic_vector(0 downto 0);
  signal readVector_call_acks: std_logic_vector(0 downto 0);
  signal readVector_return_reqs: std_logic_vector(0 downto 0);
  signal readVector_return_acks: std_logic_vector(0 downto 0);
  signal readVector_call_tag: std_logic_vector(0 downto 0);
  signal readVector_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendVector
  component sendVector is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(4 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendVector
  signal sendVector_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendVector_tag_out   : std_logic_vector(1 downto 0);
  signal sendVector_start_req : std_logic;
  signal sendVector_start_ack : std_logic;
  signal sendVector_fin_req   : std_logic;
  signal sendVector_fin_ack : std_logic;
  -- caller side aggregated signals for module sendVector
  signal sendVector_call_reqs: std_logic_vector(0 downto 0);
  signal sendVector_call_acks: std_logic_vector(0 downto 0);
  signal sendVector_return_reqs: std_logic_vector(0 downto 0);
  signal sendVector_return_acks: std_logic_vector(0 downto 0);
  signal sendVector_call_tag: std_logic_vector(0 downto 0);
  signal sendVector_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(1 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module dotP_even
  dotP_even_R <= dotP_even_in_args(7 downto 0);
  dotP_even_out_args <= dotP_even_result ;
  -- call arbiter for module dotP_even
  dotP_even_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 8,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => dotP_even_call_reqs,
      call_acks => dotP_even_call_acks,
      return_reqs => dotP_even_return_reqs,
      return_acks => dotP_even_return_acks,
      call_data  => dotP_even_call_data,
      call_tag  => dotP_even_call_tag,
      return_tag  => dotP_even_return_tag,
      call_mtag => dotP_even_tag_in,
      return_mtag => dotP_even_tag_out,
      return_data =>dotP_even_return_data,
      call_mreq => dotP_even_start_req,
      call_mack => dotP_even_start_ack,
      return_mreq => dotP_even_fin_req,
      return_mack => dotP_even_fin_ack,
      call_mdata => dotP_even_in_args,
      return_mdata => dotP_even_out_args,
      clk => clk, 
      reset => reset --
    ); --
  dotP_even_instance:dotP_even-- 
    generic map(tag_length => 2)
    port map(-- 
      R => dotP_even_R,
      result => dotP_even_result,
      start_req => dotP_even_start_req,
      start_ack => dotP_even_start_ack,
      fin_req => dotP_even_fin_req,
      fin_ack => dotP_even_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(15 downto 8),
      memory_space_0_lr_tag => memory_space_0_lr_tag(35 downto 18),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(15 downto 8),
      memory_space_1_lr_tag => memory_space_1_lr_tag(35 downto 18),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(15 downto 8),
      memory_space_2_lr_tag => memory_space_2_lr_tag(35 downto 18),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 1),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(15 downto 8),
      memory_space_3_lr_tag => memory_space_3_lr_tag(35 downto 18),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 1),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(5 downto 3),
      memory_space_4_lr_tag => memory_space_4_lr_tag(35 downto 18),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 32),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 1),
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(5 downto 3),
      memory_space_5_lr_tag => memory_space_5_lr_tag(35 downto 18),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(1 downto 1),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(5 downto 3),
      memory_space_6_lr_tag => memory_space_6_lr_tag(35 downto 18),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(5 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(35 downto 18),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 1),
      tag_in => dotP_even_tag_in,
      tag_out => dotP_even_tag_out-- 
    ); -- 
  -- module dotP_odd
  dotP_odd_R <= dotP_odd_in_args(7 downto 0);
  dotP_odd_out_args <= dotP_odd_result ;
  -- call arbiter for module dotP_odd
  dotP_odd_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 8,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => dotP_odd_call_reqs,
      call_acks => dotP_odd_call_acks,
      return_reqs => dotP_odd_return_reqs,
      return_acks => dotP_odd_return_acks,
      call_data  => dotP_odd_call_data,
      call_tag  => dotP_odd_call_tag,
      return_tag  => dotP_odd_return_tag,
      call_mtag => dotP_odd_tag_in,
      return_mtag => dotP_odd_tag_out,
      return_data =>dotP_odd_return_data,
      call_mreq => dotP_odd_start_req,
      call_mack => dotP_odd_start_ack,
      return_mreq => dotP_odd_fin_req,
      return_mack => dotP_odd_fin_ack,
      call_mdata => dotP_odd_in_args,
      return_mdata => dotP_odd_out_args,
      clk => clk, 
      reset => reset --
    ); --
  dotP_odd_instance:dotP_odd-- 
    generic map(tag_length => 2)
    port map(-- 
      R => dotP_odd_R,
      result => dotP_odd_result,
      start_req => dotP_odd_start_req,
      start_ack => dotP_odd_start_ack,
      fin_req => dotP_odd_fin_req,
      fin_ack => dotP_odd_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(7 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(7 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(7 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(7 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(17 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(2 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(17 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(2 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(17 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(17 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(17 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      tag_in => dotP_odd_tag_in,
      tag_out => dotP_odd_tag_out-- 
    ); -- 
  -- module multiplyMatrixVector
  -- call arbiter for module multiplyMatrixVector
  multiplyMatrixVector_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => multiplyMatrixVector_call_reqs,
      call_acks => multiplyMatrixVector_call_acks,
      return_reqs => multiplyMatrixVector_return_reqs,
      return_acks => multiplyMatrixVector_return_acks,
      call_tag  => multiplyMatrixVector_call_tag,
      return_tag  => multiplyMatrixVector_return_tag,
      call_mtag => multiplyMatrixVector_tag_in,
      return_mtag => multiplyMatrixVector_tag_out,
      call_mreq => multiplyMatrixVector_start_req,
      call_mack => multiplyMatrixVector_start_ack,
      return_mreq => multiplyMatrixVector_fin_req,
      return_mack => multiplyMatrixVector_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  multiplyMatrixVector_instance:multiplyMatrixVector-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => multiplyMatrixVector_start_req,
      start_ack => multiplyMatrixVector_start_ack,
      fin_req => multiplyMatrixVector_fin_req,
      fin_ack => multiplyMatrixVector_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(4 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(31 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(18 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(1 downto 0),
      dotP_even_call_reqs => dotP_even_call_reqs(0 downto 0),
      dotP_even_call_acks => dotP_even_call_acks(0 downto 0),
      dotP_even_call_data => dotP_even_call_data(7 downto 0),
      dotP_even_call_tag => dotP_even_call_tag(0 downto 0),
      dotP_even_return_reqs => dotP_even_return_reqs(0 downto 0),
      dotP_even_return_acks => dotP_even_return_acks(0 downto 0),
      dotP_even_return_data => dotP_even_return_data(31 downto 0),
      dotP_even_return_tag => dotP_even_return_tag(0 downto 0),
      dotP_odd_call_reqs => dotP_odd_call_reqs(0 downto 0),
      dotP_odd_call_acks => dotP_odd_call_acks(0 downto 0),
      dotP_odd_call_data => dotP_odd_call_data(7 downto 0),
      dotP_odd_call_tag => dotP_odd_call_tag(0 downto 0),
      dotP_odd_return_reqs => dotP_odd_return_reqs(0 downto 0),
      dotP_odd_return_acks => dotP_odd_return_acks(0 downto 0),
      dotP_odd_return_data => dotP_odd_return_data(31 downto 0),
      dotP_odd_return_tag => dotP_odd_return_tag(0 downto 0),
      tag_in => multiplyMatrixVector_tag_in,
      tag_out => multiplyMatrixVector_tag_out-- 
    ); -- 
  -- module mvp_daemon
  mvp_daemon_instance:mvp_daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => mvp_daemon_start_req,
      start_ack => mvp_daemon_start_ack,
      fin_req => mvp_daemon_fin_req,
      fin_ack => mvp_daemon_fin_ack,
      clk => clk,
      reset => reset,
      multiplyMatrixVector_call_reqs => multiplyMatrixVector_call_reqs(0 downto 0),
      multiplyMatrixVector_call_acks => multiplyMatrixVector_call_acks(0 downto 0),
      multiplyMatrixVector_call_tag => multiplyMatrixVector_call_tag(0 downto 0),
      multiplyMatrixVector_return_reqs => multiplyMatrixVector_return_reqs(0 downto 0),
      multiplyMatrixVector_return_acks => multiplyMatrixVector_return_acks(0 downto 0),
      multiplyMatrixVector_return_tag => multiplyMatrixVector_return_tag(0 downto 0),
      readMatrix_call_reqs => readMatrix_call_reqs(0 downto 0),
      readMatrix_call_acks => readMatrix_call_acks(0 downto 0),
      readMatrix_call_tag => readMatrix_call_tag(0 downto 0),
      readMatrix_return_reqs => readMatrix_return_reqs(0 downto 0),
      readMatrix_return_acks => readMatrix_return_acks(0 downto 0),
      readMatrix_return_tag => readMatrix_return_tag(0 downto 0),
      readVector_call_reqs => readVector_call_reqs(0 downto 0),
      readVector_call_acks => readVector_call_acks(0 downto 0),
      readVector_call_tag => readVector_call_tag(0 downto 0),
      readVector_return_reqs => readVector_return_reqs(0 downto 0),
      readVector_return_acks => readVector_return_acks(0 downto 0),
      readVector_return_tag => readVector_return_tag(0 downto 0),
      sendVector_call_reqs => sendVector_call_reqs(0 downto 0),
      sendVector_call_acks => sendVector_call_acks(0 downto 0),
      sendVector_call_tag => sendVector_call_tag(0 downto 0),
      sendVector_return_reqs => sendVector_return_reqs(0 downto 0),
      sendVector_return_acks => sendVector_return_acks(0 downto 0),
      sendVector_return_tag => sendVector_return_tag(0 downto 0),
      tag_in => mvp_daemon_tag_in,
      tag_out => mvp_daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  mvp_daemon_tag_in <= (others => '0');
  mvp_daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => mvp_daemon_start_req, start_ack => mvp_daemon_start_ack,  fin_req => mvp_daemon_fin_req,  fin_ack => mvp_daemon_fin_ack);
  -- module readMatrix
  -- call arbiter for module readMatrix
  readMatrix_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readMatrix_call_reqs,
      call_acks => readMatrix_call_acks,
      return_reqs => readMatrix_return_reqs,
      return_acks => readMatrix_return_acks,
      call_tag  => readMatrix_call_tag,
      return_tag  => readMatrix_return_tag,
      call_mtag => readMatrix_tag_in,
      return_mtag => readMatrix_tag_out,
      call_mreq => readMatrix_start_req,
      call_mack => readMatrix_start_ack,
      return_mreq => readMatrix_fin_req,
      return_mack => readMatrix_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  readMatrix_instance:readMatrix-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => readMatrix_start_req,
      start_ack => readMatrix_start_ack,
      fin_req => readMatrix_fin_req,
      fin_ack => readMatrix_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(7 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(7 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(7 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(7 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(17 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(31 downto 0),
      tag_in => readMatrix_tag_in,
      tag_out => readMatrix_tag_out-- 
    ); -- 
  -- module readVector
  -- call arbiter for module readVector
  readVector_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readVector_call_reqs,
      call_acks => readVector_call_acks,
      return_reqs => readVector_return_reqs,
      return_acks => readVector_return_acks,
      call_tag  => readVector_call_tag,
      return_tag  => readVector_return_tag,
      call_mtag => readVector_tag_in,
      return_mtag => readVector_tag_out,
      call_mreq => readVector_start_req,
      call_mack => readVector_start_ack,
      return_mreq => readVector_fin_req,
      return_mack => readVector_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  readVector_instance:readVector-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => readVector_start_req,
      start_ack => readVector_start_ack,
      fin_req => readVector_fin_req,
      fin_ack => readVector_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(2 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(17 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(2 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(17 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(2 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(31 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(17 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(2 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(31 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(17 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(1 downto 1),
      in_data_pipe_read_ack => in_data_pipe_read_ack(1 downto 1),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 32),
      tag_in => readVector_tag_in,
      tag_out => readVector_tag_out-- 
    ); -- 
  -- module sendVector
  -- call arbiter for module sendVector
  sendVector_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendVector_call_reqs,
      call_acks => sendVector_call_acks,
      return_reqs => sendVector_return_reqs,
      return_acks => sendVector_return_acks,
      call_tag  => sendVector_call_tag,
      return_tag  => sendVector_return_tag,
      call_mtag => sendVector_tag_in,
      return_mtag => sendVector_tag_out,
      call_mreq => sendVector_start_req,
      call_mack => sendVector_start_ack,
      return_mreq => sendVector_fin_req,
      return_mack => sendVector_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendVector_instance:sendVector-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendVector_start_req,
      start_ack => sendVector_start_ack,
      fin_req => sendVector_fin_req,
      fin_ack => sendVector_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(4 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(18 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(1 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(31 downto 0),
      tag_in => sendVector_tag_in,
      tag_out => sendVector_tag_out-- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data",
      num_reads => 2,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 2,
      num_stores => 1,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 2,
      num_stores => 1,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 2,
      num_stores => 1,
      addr_width => 8,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 8,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 2,
      num_stores => 1,
      addr_width => 3,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 2,
      num_stores => 1,
      addr_width => 3,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 2,
      num_stores => 1,
      addr_width => 3,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 2,
      num_stores => 1,
      addr_width => 3,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 1,
      num_stores => 1,
      addr_width => 5,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 5,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;

-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant A_0_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant A_1_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant x_0_base_address : std_logic_vector(3 downto 0) := "0000";
  constant x_1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant y_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package ahir_system_global_package;
